module small_circle (
    input wire Gi,
    output wire Ci
);
  
  assign Ci = Gi;
  
endmodule