
`timescale 1ns / 1ps

module tb_N7_booth_multiplier;

    // Parameters
    
    parameter N = 7;
    
     
    // Inputs
    
    reg   clk;
    
    reg   rst;
    
    reg   start;
    
    reg signed [6:0] X;
    
    reg signed [6:0] Y;
    
    
    // Outputs
    
    wire signed [13:0] Z;
    
    wire   valid;
    
    
    // Instantiate the Unit Under Test (UUT)
    booth_multiplier  #( N ) uut (
        
        .clk(clk),
        
        .rst(rst),
        
        .start(start),
        
        .X(X),
        
        .Y(Y),
        
        
        .Z(Z),
        
        .valid(valid)
        
    );

    // Clock generation 
    
    
            always begin
                #5 clk = ~clk;
            end
            
    

    
    
            always begin
                #99 rst = 1'b1; 
            end
            
    
    
    initial begin
        // Initialize Inputs
        
        clk = 0;
        
        rst = 0;
        
        start = 0;
        
        X = 0;
        
        Y = 0;
        
    
        // Wait for global reset
        #100;
    
        // Stimuli
        
        #10 X = 7'b1000000; Y = 7'b1011100; // Expected: {'Z': 2304}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000000; Y = 7'b1011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 0,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2304
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111010; Y = 7'b1101001; // Expected: {'Z': 138}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111010; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011111; Y = 7'b1100000; // Expected: {'Z': -992}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011111; Y = 7'b1100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -992
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b0101011; // Expected: {'Z': 43}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b0101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101000; Y = 7'b0110000; // Expected: {'Z': 1920}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101000; Y = 7'b0110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 4,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b1011111; // Expected: {'Z': -1485}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 5,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1485
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100001; Y = 7'b0111100; // Expected: {'Z': 1980}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100001; Y = 7'b0111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 6,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b0100111; // Expected: {'Z': 1755}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b0100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 7,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1755
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100001; Y = 7'b0010000; // Expected: {'Z': 528}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100001; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 8,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101111; Y = 7'b0001000; // Expected: {'Z': 376}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101111; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 9,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 376
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b0010110; // Expected: {'Z': -22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b0010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 10,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110000; Y = 7'b1100011; // Expected: {'Z': -1392}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110000; Y = 7'b1100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 11,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b1010001; // Expected: {'Z': 2961}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 12,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2961
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100000; Y = 7'b0011010; // Expected: {'Z': 832}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100000; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 13,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 832
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b1011000; // Expected: {'Z': 1120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b1011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 14,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b1110101; // Expected: {'Z': 440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b1110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 15,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110101; Y = 7'b0011000; // Expected: {'Z': -264}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110101; Y = 7'b0011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 16,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001000; Y = 7'b1010100; // Expected: {'Z': -352}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001000; Y = 7'b1010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 17,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100001; Y = 7'b0000100; // Expected: {'Z': 132}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100001; Y = 7'b0000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 18,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100011; Y = 7'b0110101; // Expected: {'Z': -1537}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100011; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 19,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1537
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010010; Y = 7'b0001111; // Expected: {'Z': 270}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010010; Y = 7'b0001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 20,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 270
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111010; Y = 7'b0111001; // Expected: {'Z': -342}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111010; Y = 7'b0111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 21,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -342
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b1100111; // Expected: {'Z': 75}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b1100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 22,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b1000100; // Expected: {'Z': 900}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b1000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 23,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110111; Y = 7'b1000110; // Expected: {'Z': 522}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110111; Y = 7'b1000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 24,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 522
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b0101111; // Expected: {'Z': 940}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b0101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 25,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 940
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001100; Y = 7'b0100101; // Expected: {'Z': 444}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001100; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 26,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 444
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b0010001; // Expected: {'Z': -51}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 27,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010100; Y = 7'b1101100; // Expected: {'Z': 880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010100; Y = 7'b1101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 28,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b1001001; // Expected: {'Z': 2640}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b1001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 29,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000111; Y = 7'b0001001; // Expected: {'Z': 63}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000111; Y = 7'b0001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 30,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110111; Y = 7'b1101100; // Expected: {'Z': 180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110111; Y = 7'b1101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 31,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110001; Y = 7'b0011110; // Expected: {'Z': 1470}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110001; Y = 7'b0011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 32,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1470
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110010; Y = 7'b0110010; // Expected: {'Z': -700}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110010; Y = 7'b0110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 33,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100111; Y = 7'b0110000; // Expected: {'Z': 1872}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100111; Y = 7'b0110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 34,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1872
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110110; Y = 7'b0100010; // Expected: {'Z': 1836}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110110; Y = 7'b0100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 35,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1836
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101000; Y = 7'b1110010; // Expected: {'Z': -560}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101000; Y = 7'b1110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 36,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000010; Y = 7'b1001011; // Expected: {'Z': 3286}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000010; Y = 7'b1001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 37,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3286
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100111; Y = 7'b1110111; // Expected: {'Z': -351}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100111; Y = 7'b1110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 38,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -351
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100111; Y = 7'b0011000; // Expected: {'Z': -600}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100111; Y = 7'b0011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 39,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000111; Y = 7'b1001111; // Expected: {'Z': -343}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000111; Y = 7'b1001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 40,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -343
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011101; Y = 7'b0100010; // Expected: {'Z': -1190}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011101; Y = 7'b0100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 41,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011110; Y = 7'b0000111; // Expected: {'Z': 210}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011110; Y = 7'b0000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 42,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101011; Y = 7'b0011001; // Expected: {'Z': -525}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101011; Y = 7'b0011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 43,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -525
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101110; Y = 7'b0111101; // Expected: {'Z': 2806}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101110; Y = 7'b0111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 44,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2806
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011101; Y = 7'b0010111; // Expected: {'Z': 667}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011101; Y = 7'b0010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 45,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 667
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110011; Y = 7'b0101010; // Expected: {'Z': 2142}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110011; Y = 7'b0101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 46,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010001; Y = 7'b1111101; // Expected: {'Z': 141}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010001; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 47,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101011; Y = 7'b1010011; // Expected: {'Z': -1935}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101011; Y = 7'b1010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 48,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1935
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b1100101; // Expected: {'Z': -648}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 49,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000010; Y = 7'b1110000; // Expected: {'Z': 992}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000010; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 50,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 992
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100000; Y = 7'b1010000; // Expected: {'Z': -1536}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100000; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 51,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1536
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b0111010; // Expected: {'Z': 58}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 52,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b1111100; // Expected: {'Z': 128}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 53,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b0110101; // Expected: {'Z': -1060}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 54,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b1001110; // Expected: {'Z': -1000}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b1001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 55,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101011; Y = 7'b0010001; // Expected: {'Z': -357}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101011; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 56,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -357
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b1111001; // Expected: {'Z': 441}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b1111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 57,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 441
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b1010011; // Expected: {'Z': 765}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b1010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 58,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 765
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111010; Y = 7'b0110110; // Expected: {'Z': -324}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111010; Y = 7'b0110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 59,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -324
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111010; Y = 7'b1101111; // Expected: {'Z': -986}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111010; Y = 7'b1101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 60,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -986
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010010; Y = 7'b0011100; // Expected: {'Z': 504}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010010; Y = 7'b0011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 61,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b1111100; // Expected: {'Z': 80}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 62,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110111; Y = 7'b1111111; // Expected: {'Z': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110111; Y = 7'b1111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 63,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110010; Y = 7'b1000000; // Expected: {'Z': 896}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110010; Y = 7'b1000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 64,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001010; Y = 7'b0101001; // Expected: {'Z': 410}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001010; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 65,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 410
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b1100011; // Expected: {'Z': 1392}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b1100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 66,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111001; Y = 7'b1000011; // Expected: {'Z': -3477}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111001; Y = 7'b1000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 67,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3477
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000010; Y = 7'b0001001; // Expected: {'Z': -558}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000010; Y = 7'b0001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 68,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -558
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b1111001; // Expected: {'Z': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b1111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 69,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001000; Y = 7'b1100000; // Expected: {'Z': -256}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001000; Y = 7'b1100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 70,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -256
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111010; Y = 7'b0000111; // Expected: {'Z': 406}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111010; Y = 7'b0000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 71,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 406
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110010; Y = 7'b0101001; // Expected: {'Z': 2050}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110010; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 72,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b1100010; // Expected: {'Z': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 73,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000101; Y = 7'b0100010; // Expected: {'Z': -2006}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000101; Y = 7'b0100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 74,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2006
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010000; Y = 7'b1001011; // Expected: {'Z': -848}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010000; Y = 7'b1001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 75,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111001; Y = 7'b1101011; // Expected: {'Z': -1197}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111001; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 76,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011101; Y = 7'b0001000; // Expected: {'Z': -280}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011101; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 77,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101110; Y = 7'b1100100; // Expected: {'Z': -1288}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101110; Y = 7'b1100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 78,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010111; Y = 7'b0101001; // Expected: {'Z': 943}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010111; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 79,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 943
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100100; Y = 7'b0110111; // Expected: {'Z': 1980}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100100; Y = 7'b0110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 80,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010110; Y = 7'b1101011; // Expected: {'Z': -462}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010110; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 81,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110010; Y = 7'b1011111; // Expected: {'Z': 462}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110010; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 82,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011011; Y = 7'b0111010; // Expected: {'Z': -2146}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011011; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 83,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100001; Y = 7'b0001111; // Expected: {'Z': 495}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100001; Y = 7'b0001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 84,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 495
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000000; Y = 7'b1000010; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000000; Y = 7'b1000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 85,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011001; Y = 7'b0101100; // Expected: {'Z': 1100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011001; Y = 7'b0101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 86,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100110; Y = 7'b0010000; // Expected: {'Z': 608}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100110; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 87,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 608
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b1100010; // Expected: {'Z': 1200}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 88,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b1111001; // Expected: {'Z': -147}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b1111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 89,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111000; Y = 7'b0010000; // Expected: {'Z': 896}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111000; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 90,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100010; Y = 7'b1101011; // Expected: {'Z': -714}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100010; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 91,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -714
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011110; Y = 7'b1110000; // Expected: {'Z': -480}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011110; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 92,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b1001001; // Expected: {'Z': -2915}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b1001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 93,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2915
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001001; Y = 7'b0010110; // Expected: {'Z': -1210}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001001; Y = 7'b0010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 94,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010010; Y = 7'b1111011; // Expected: {'Z': 230}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010010; Y = 7'b1111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 95,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101011; Y = 7'b1001110; // Expected: {'Z': -2150}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101011; Y = 7'b1001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 96,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011001; Y = 7'b0111001; // Expected: {'Z': -2223}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011001; Y = 7'b0111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 97,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2223
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110011; Y = 7'b0010011; // Expected: {'Z': -247}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110011; Y = 7'b0010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 98,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001000; Y = 7'b0100101; // Expected: {'Z': 296}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001000; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 99,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001110; Y = 7'b0010011; // Expected: {'Z': -950}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001110; Y = 7'b0010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 100,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101000; Y = 7'b1110001; // Expected: {'Z': -600}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101000; Y = 7'b1110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 101,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b1101001; // Expected: {'Z': 1449}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 102,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1449
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101010; Y = 7'b1000111; // Expected: {'Z': -2394}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101010; Y = 7'b1000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 103,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2394
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b0110010; // Expected: {'Z': -900}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b0110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 104,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000000; Y = 7'b0100001; // Expected: {'Z': -2112}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000000; Y = 7'b0100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 105,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111000; Y = 7'b0001101; // Expected: {'Z': -104}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111000; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 106,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011100; Y = 7'b1000100; // Expected: {'Z': -1680}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011100; Y = 7'b1000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 107,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000100; Y = 7'b1000000; // Expected: {'Z': -256}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000100; Y = 7'b1000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 108,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -256
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b0111010; // Expected: {'Z': -2088}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 109,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2088
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110111; Y = 7'b0111011; // Expected: {'Z': 3245}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110111; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 110,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100010; Y = 7'b0001000; // Expected: {'Z': 272}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100010; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 111,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 272
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100100; Y = 7'b1011001; // Expected: {'Z': -1404}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100100; Y = 7'b1011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 112,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1404
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111001; Y = 7'b1001000; // Expected: {'Z': -3192}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111001; Y = 7'b1001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 113,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b0001001; // Expected: {'Z': 180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b0001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 114,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000010; Y = 7'b0010010; // Expected: {'Z': -1116}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000010; Y = 7'b0010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 115,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100111; Y = 7'b1000010; // Expected: {'Z': -2418}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100111; Y = 7'b1000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 116,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2418
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111001; Y = 7'b0000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111001; Y = 7'b0000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 117,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100111; Y = 7'b0100010; // Expected: {'Z': -850}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100111; Y = 7'b0100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 118,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -850
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100111; Y = 7'b0100100; // Expected: {'Z': 1404}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100111; Y = 7'b0100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 119,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1404
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100001; Y = 7'b1010010; // Expected: {'Z': -1518}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100001; Y = 7'b1010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 120,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1518
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001110; Y = 7'b0100011; // Expected: {'Z': -1750}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001110; Y = 7'b0100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 121,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b1101101; // Expected: {'Z': 323}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b1101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 122,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 323
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b0011100; // Expected: {'Z': -1764}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b0011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 123,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1764
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110111; Y = 7'b1110011; // Expected: {'Z': -715}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110111; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 124,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -715
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b1101111; // Expected: {'Z': 680}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b1101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 125,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000111; Y = 7'b1001101; // Expected: {'Z': -357}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000111; Y = 7'b1001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 126,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -357
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b1111011; // Expected: {'Z': 140}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b1111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 127,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b0111001; // Expected: {'Z': -1938}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b0111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 128,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1938
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101010; Y = 7'b1010110; // Expected: {'Z': 924}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101010; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 129,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 924
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000110; Y = 7'b1101001; // Expected: {'Z': 1334}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000110; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 130,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1334
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b1001000; // Expected: {'Z': 952}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b1001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 131,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 952
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000100; Y = 7'b1011011; // Expected: {'Z': 2220}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000100; Y = 7'b1011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 132,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000010; Y = 7'b0110100; // Expected: {'Z': 104}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000010; Y = 7'b0110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 133,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110010; Y = 7'b0101100; // Expected: {'Z': -616}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110010; Y = 7'b0101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 134,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -616
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101010; Y = 7'b0110110; // Expected: {'Z': 2268}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101010; Y = 7'b0110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 135,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2268
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010101; Y = 7'b0100111; // Expected: {'Z': -1677}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010101; Y = 7'b0100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 136,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1677
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b0100110; // Expected: {'Z': 2356}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 137,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2356
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111001; Y = 7'b1010111; // Expected: {'Z': -2337}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111001; Y = 7'b1010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 138,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2337
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b1011001; // Expected: {'Z': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b1011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 139,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101010; Y = 7'b0000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101010; Y = 7'b0000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 140,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001100; Y = 7'b0111010; // Expected: {'Z': -3016}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001100; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 141,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101000; Y = 7'b0111011; // Expected: {'Z': -1416}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101000; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 142,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011011; Y = 7'b0100000; // Expected: {'Z': -1184}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011011; Y = 7'b0100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 143,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b1010000; // Expected: {'Z': 48}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 144,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000101; Y = 7'b0100100; // Expected: {'Z': 180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000101; Y = 7'b0100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 145,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b1100001; // Expected: {'Z': 465}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b1100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 146,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 465
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b1011100; // Expected: {'Z': -1620}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b1011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 147,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011101; Y = 7'b0010111; // Expected: {'Z': -805}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011101; Y = 7'b0010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 148,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -805
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000111; Y = 7'b1110100; // Expected: {'Z': -84}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000111; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 149,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b1101101; // Expected: {'Z': 228}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b1101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 150,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001111; Y = 7'b1110100; // Expected: {'Z': -180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001111; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 151,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001100; Y = 7'b0000100; // Expected: {'Z': -208}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001100; Y = 7'b0000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 152,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b0100101; // Expected: {'Z': -666}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 153,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -666
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001100; Y = 7'b1001010; // Expected: {'Z': 2808}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001100; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 154,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001010; Y = 7'b1010000; // Expected: {'Z': 2592}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001010; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 155,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2592
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001110; Y = 7'b1111111; // Expected: {'Z': -14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001110; Y = 7'b1111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 156,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b0101011; // Expected: {'Z': -1720}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b0101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 157,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001000; Y = 7'b1101001; // Expected: {'Z': -184}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001000; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 158,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010000; Y = 7'b1000011; // Expected: {'Z': -976}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010000; Y = 7'b1000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 159,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -976
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111110; Y = 7'b0110100; // Expected: {'Z': -104}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111110; Y = 7'b0110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 160,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010101; Y = 7'b1101110; // Expected: {'Z': 774}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010101; Y = 7'b1101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 161,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 774
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b1001000; // Expected: {'Z': 1792}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b1001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 162,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010010; Y = 7'b0111010; // Expected: {'Z': 1044}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010010; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 163,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1044
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111100; Y = 7'b1100101; // Expected: {'Z': 108}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111100; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 164,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011011; Y = 7'b0100101; // Expected: {'Z': 999}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011011; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 165,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 999
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000010; Y = 7'b0111110; // Expected: {'Z': -3844}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000010; Y = 7'b0111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 166,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3844
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010001; Y = 7'b0101100; // Expected: {'Z': -2068}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010001; Y = 7'b0101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 167,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2068
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101011; Y = 7'b1011010; // Expected: {'Z': -1634}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101011; Y = 7'b1011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 168,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1634
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100011; Y = 7'b1011101; // Expected: {'Z': -1225}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100011; Y = 7'b1011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 169,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101110; Y = 7'b0101100; // Expected: {'Z': 2024}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101110; Y = 7'b0101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 170,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b0001101; // Expected: {'Z': 585}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 171,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 585
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101010; Y = 7'b1011010; // Expected: {'Z': -1596}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101010; Y = 7'b1011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 172,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1596
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001001; Y = 7'b1110110; // Expected: {'Z': 550}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001001; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 173,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101011; Y = 7'b1001010; // Expected: {'Z': -2322}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101011; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 174,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2322
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001110; Y = 7'b0011000; // Expected: {'Z': -1200}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001110; Y = 7'b0011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 175,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b0001011; // Expected: {'Z': 187}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b0001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 176,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000101; Y = 7'b0100001; // Expected: {'Z': 165}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000101; Y = 7'b0100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 177,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001000; Y = 7'b0000010; // Expected: {'Z': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001000; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 178,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b0100000; // Expected: {'Z': -384}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b0100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 179,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -384
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110110; Y = 7'b0111000; // Expected: {'Z': 3024}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110110; Y = 7'b0111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 180,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110001; Y = 7'b0110111; // Expected: {'Z': 2695}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110001; Y = 7'b0110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 181,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2695
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111001; Y = 7'b1111100; // Expected: {'Z': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111001; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 182,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b1111110; // Expected: {'Z': 40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b1111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 183,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101000; Y = 7'b0101001; // Expected: {'Z': 1640}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101000; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 184,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011011; Y = 7'b1000011; // Expected: {'Z': -1647}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011011; Y = 7'b1000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 185,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1647
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b0001110; // Expected: {'Z': -588}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 186,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -588
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111111; Y = 7'b0111010; // Expected: {'Z': 3654}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111111; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 187,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3654
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b0000010; // Expected: {'Z': -6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 188,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011111; Y = 7'b0010011; // Expected: {'Z': 589}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011111; Y = 7'b0010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 189,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 589
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111101; Y = 7'b1110110; // Expected: {'Z': -610}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111101; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 190,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -610
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b0010000; // Expected: {'Z': -160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 191,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100111; Y = 7'b0010010; // Expected: {'Z': 702}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100111; Y = 7'b0010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 192,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 702
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010010; Y = 7'b0100110; // Expected: {'Z': -1748}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010010; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 193,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1748
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011110; Y = 7'b1001110; // Expected: {'Z': -1500}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011110; Y = 7'b1001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 194,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b0000111; // Expected: {'Z': -294}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b0000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 195,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -294
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011001; Y = 7'b1101100; // Expected: {'Z': -500}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011001; Y = 7'b1101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 196,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100101; Y = 7'b1101001; // Expected: {'Z': 621}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100101; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 197,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 621
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111110; Y = 7'b1111100; // Expected: {'Z': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111110; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 198,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b1010011; // Expected: {'Z': -135}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b1010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 199,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011010; Y = 7'b0100111; // Expected: {'Z': 1014}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011010; Y = 7'b0100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 200,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1014
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110001; Y = 7'b0011011; // Expected: {'Z': 1323}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110001; Y = 7'b0011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 201,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1323
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100101; Y = 7'b0010010; // Expected: {'Z': -486}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100101; Y = 7'b0010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 202,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -486
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011101; Y = 7'b1100101; // Expected: {'Z': 945}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011101; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 203,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 945
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110011; Y = 7'b1011101; // Expected: {'Z': 455}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110011; Y = 7'b1011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 204,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 455
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011010; Y = 7'b1111111; // Expected: {'Z': -26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011010; Y = 7'b1111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 205,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b0111101; // Expected: {'Z': -1403}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b0111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 206,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1403
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b1101111; // Expected: {'Z': 306}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b1101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 207,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 306
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101111; Y = 7'b0000110; // Expected: {'Z': 282}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101111; Y = 7'b0000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 208,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 282
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110000; Y = 7'b1011011; // Expected: {'Z': -1776}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110000; Y = 7'b1011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 209,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1776
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110011; Y = 7'b0100101; // Expected: {'Z': 1887}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110011; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 210,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1887
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010111; Y = 7'b1111000; // Expected: {'Z': -184}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010111; Y = 7'b1111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 211,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b0010001; // Expected: {'Z': 51}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 212,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110111; Y = 7'b0101111; // Expected: {'Z': -423}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110111; Y = 7'b0101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 213,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -423
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110000; Y = 7'b1110100; // Expected: {'Z': 192}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110000; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 214,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011111; Y = 7'b0101001; // Expected: {'Z': -1353}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011111; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 215,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1353
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b0100100; // Expected: {'Z': -1008}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b0100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 216,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b1010111; // Expected: {'Z': 492}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b1010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 217,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 492
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001101; Y = 7'b0110011; // Expected: {'Z': -2601}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001101; Y = 7'b0110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 218,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2601
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b0101011; // Expected: {'Z': 2666}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b0101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 219,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2666
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111001; Y = 7'b1011000; // Expected: {'Z': 280}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111001; Y = 7'b1011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 220,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010100; Y = 7'b0100101; // Expected: {'Z': -1628}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010100; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 221,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1628
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111010; Y = 7'b0000101; // Expected: {'Z': -30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111010; Y = 7'b0000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 222,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110010; Y = 7'b1101100; // Expected: {'Z': 280}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110010; Y = 7'b1101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 223,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101110; Y = 7'b0011111; // Expected: {'Z': 1426}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101110; Y = 7'b0011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 224,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1426
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b0011001; // Expected: {'Z': -1200}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b0011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 225,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011011; Y = 7'b0010100; // Expected: {'Z': 540}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011011; Y = 7'b0010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 226,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011010; Y = 7'b0100111; // Expected: {'Z': -1482}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011010; Y = 7'b0100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 227,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1482
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b1111110; // Expected: {'Z': 34}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b1111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 228,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001001; Y = 7'b0011000; // Expected: {'Z': -1320}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001001; Y = 7'b0011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 229,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b1111100; // Expected: {'Z': -248}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 230,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001100; Y = 7'b1110010; // Expected: {'Z': 728}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001100; Y = 7'b1110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 231,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011001; Y = 7'b1001000; // Expected: {'Z': -1400}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011001; Y = 7'b1001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 232,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100111; Y = 7'b1000111; // Expected: {'Z': 1425}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100111; Y = 7'b1000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 233,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1425
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b0000001; // Expected: {'Z': 45}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b0000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 234,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000010; Y = 7'b0001110; // Expected: {'Z': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000010; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 235,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b0010110; // Expected: {'Z': 66}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b0010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 236,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b0100011; // Expected: {'Z': 2170}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b0100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 237,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101001; Y = 7'b1101000; // Expected: {'Z': -984}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101001; Y = 7'b1101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 238,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -984
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010110; Y = 7'b1010000; // Expected: {'Z': -1056}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010110; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 239,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1056
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000100; Y = 7'b1101001; // Expected: {'Z': -92}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000100; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 240,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b0100001; // Expected: {'Z': -99}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b0100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 241,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b1100110; // Expected: {'Z': -546}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b1100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 242,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110110; Y = 7'b0001100; // Expected: {'Z': 648}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110110; Y = 7'b0001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 243,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101111; Y = 7'b0111011; // Expected: {'Z': 2773}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101111; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 244,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2773
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010000; Y = 7'b1100000; // Expected: {'Z': -512}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010000; Y = 7'b1100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 245,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -512
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111000; Y = 7'b1010111; // Expected: {'Z': 328}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111000; Y = 7'b1010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 246,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 328
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101110; Y = 7'b0101001; // Expected: {'Z': 1886}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101110; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 247,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1886
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101001; Y = 7'b1001101; // Expected: {'Z': -2091}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101001; Y = 7'b1001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 248,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2091
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101000; Y = 7'b0001001; // Expected: {'Z': 360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101000; Y = 7'b0001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 249,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100110; Y = 7'b0011101; // Expected: {'Z': 1102}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100110; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 250,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001101; Y = 7'b1000100; // Expected: {'Z': -780}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001101; Y = 7'b1000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 251,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b1001101; // Expected: {'Z': 2142}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b1001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 252,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001101; Y = 7'b1101100; // Expected: {'Z': 1020}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001101; Y = 7'b1101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 253,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1020
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101110; Y = 7'b1010001; // Expected: {'Z': -2162}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101110; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 254,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110010; Y = 7'b1111001; // Expected: {'Z': -350}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110010; Y = 7'b1111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 255,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b1010000; // Expected: {'Z': 3024}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 256,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110001; Y = 7'b1101000; // Expected: {'Z': -1176}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110001; Y = 7'b1101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 257,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110111; Y = 7'b1111000; // Expected: {'Z': 72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110111; Y = 7'b1111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 258,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b1110010; // Expected: {'Z': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b1110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 259,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001110; Y = 7'b1100101; // Expected: {'Z': -378}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001110; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 260,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -378
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101110; Y = 7'b0110010; // Expected: {'Z': 2300}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101110; Y = 7'b0110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 261,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100110; Y = 7'b0000111; // Expected: {'Z': -182}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100110; Y = 7'b0000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 262,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b0110011; // Expected: {'Z': 51}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b0110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 263,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b1011010; // Expected: {'Z': -798}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b1011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 264,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000101; Y = 7'b1011101; // Expected: {'Z': 2065}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000101; Y = 7'b1011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 265,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2065
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b1010011; // Expected: {'Z': -765}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b1010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 266,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -765
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001101; Y = 7'b1110000; // Expected: {'Z': -208}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001101; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 267,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010111; Y = 7'b0011011; // Expected: {'Z': -1107}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010111; Y = 7'b0011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 268,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101010; Y = 7'b0001011; // Expected: {'Z': 462}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101010; Y = 7'b0001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 269,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101110; Y = 7'b1110111; // Expected: {'Z': -414}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101110; Y = 7'b1110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 270,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -414
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b1000000; // Expected: {'Z': -1280}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b1000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 271,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b1100001; // Expected: {'Z': -527}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b1100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 272,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -527
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100110; Y = 7'b0111001; // Expected: {'Z': 2166}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100110; Y = 7'b0111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 273,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001111; Y = 7'b0111101; // Expected: {'Z': -2989}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001111; Y = 7'b0111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 274,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2989
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001000; Y = 7'b1101001; // Expected: {'Z': 1288}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001000; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 275,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010111; Y = 7'b1100010; // Expected: {'Z': -690}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010111; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 276,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -690
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101011; Y = 7'b1010001; // Expected: {'Z': 987}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101011; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 277,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 987
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110011; Y = 7'b0111111; // Expected: {'Z': -819}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110011; Y = 7'b0111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 278,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -819
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b0110111; // Expected: {'Z': 495}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b0110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 279,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 495
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b0100100; // Expected: {'Z': -1728}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b0100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 280,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111011; Y = 7'b0010001; // Expected: {'Z': 1003}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111011; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 281,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1003
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b1100110; // Expected: {'Z': 494}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b1100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 282,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 494
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b1010011; // Expected: {'Z': 675}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b1010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 283,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 675
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b1101001; // Expected: {'Z': -23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 284,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b1000000; // Expected: {'Z': 1920}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b1000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 285,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010010; Y = 7'b1100111; // Expected: {'Z': -450}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010010; Y = 7'b1100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 286,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010000; Y = 7'b0011010; // Expected: {'Z': 416}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010000; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 287,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101011; Y = 7'b1000011; // Expected: {'Z': -2623}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101011; Y = 7'b1000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 288,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2623
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011011; Y = 7'b0010111; // Expected: {'Z': -851}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011011; Y = 7'b0010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 289,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -851
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110011; Y = 7'b0011111; // Expected: {'Z': 1581}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110011; Y = 7'b0011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 290,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1581
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011110; Y = 7'b0000011; // Expected: {'Z': 90}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011110; Y = 7'b0000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 291,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001011; Y = 7'b1010110; // Expected: {'Z': -462}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001011; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 292,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100100; Y = 7'b0000101; // Expected: {'Z': 180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100100; Y = 7'b0000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 293,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000100; Y = 7'b0111010; // Expected: {'Z': 232}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000100; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 294,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010101; Y = 7'b1101101; // Expected: {'Z': 817}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010101; Y = 7'b1101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 295,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 817
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b0101011; // Expected: {'Z': -430}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b0101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 296,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b0100110; // Expected: {'Z': 646}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 297,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 646
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b1111100; // Expected: {'Z': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 298,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110101; Y = 7'b1000010; // Expected: {'Z': 682}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110101; Y = 7'b1000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 299,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 682
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000100; Y = 7'b0110101; // Expected: {'Z': 212}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000100; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 300,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101010; Y = 7'b1101100; // Expected: {'Z': -840}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101010; Y = 7'b1101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 301,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001011; Y = 7'b1100000; // Expected: {'Z': -352}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001011; Y = 7'b1100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 302,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100110; Y = 7'b1011001; // Expected: {'Z': 1014}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100110; Y = 7'b1011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 303,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1014
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b1011111; // Expected: {'Z': 495}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 304,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 495
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101000; Y = 7'b1000011; // Expected: {'Z': 1464}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101000; Y = 7'b1000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 305,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b1010100; // Expected: {'Z': 880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b1010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 306,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100001; Y = 7'b1101010; // Expected: {'Z': 682}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100001; Y = 7'b1101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 307,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 682
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001110; Y = 7'b1101110; // Expected: {'Z': -252}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001110; Y = 7'b1101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 308,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b1110010; // Expected: {'Z': -630}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b1110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 309,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -630
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110000; Y = 7'b0001110; // Expected: {'Z': -224}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110000; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 310,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100001; Y = 7'b0010100; // Expected: {'Z': 660}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100001; Y = 7'b0010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 311,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b0001101; // Expected: {'Z': 117}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 312,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000100; Y = 7'b0000010; // Expected: {'Z': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000100; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 313,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000000; Y = 7'b0001011; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000000; Y = 7'b0001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 314,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011111; Y = 7'b0011110; // Expected: {'Z': -990}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011111; Y = 7'b0011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 315,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -990
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b0011010; // Expected: {'Z': 546}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 316,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011001; Y = 7'b1100110; // Expected: {'Z': 1014}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011001; Y = 7'b1100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 317,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1014
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100011; Y = 7'b0000001; // Expected: {'Z': 35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100011; Y = 7'b0000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 318,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000111; Y = 7'b1101011; // Expected: {'Z': 1197}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000111; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 319,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110101; Y = 7'b0111001; // Expected: {'Z': -627}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110101; Y = 7'b0111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 320,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -627
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b1101101; // Expected: {'Z': -19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b1101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 321,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000101; Y = 7'b1010001; // Expected: {'Z': 2773}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000101; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 322,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2773
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111011; Y = 7'b1110111; // Expected: {'Z': 45}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111011; Y = 7'b1110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 323,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100000; Y = 7'b0000110; // Expected: {'Z': 192}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100000; Y = 7'b0000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 324,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100010; Y = 7'b0100110; // Expected: {'Z': 1292}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100010; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 325,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1292
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010111; Y = 7'b1000010; // Expected: {'Z': -1426}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010111; Y = 7'b1000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 326,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1426
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101011; Y = 7'b1001001; // Expected: {'Z': -2365}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101011; Y = 7'b1001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 327,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2365
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b0101110; // Expected: {'Z': -782}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b0101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 328,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -782
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010010; Y = 7'b0000011; // Expected: {'Z': 54}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010010; Y = 7'b0000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 329,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111101; Y = 7'b0000110; // Expected: {'Z': 366}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111101; Y = 7'b0000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 330,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 366
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000110; Y = 7'b0011010; // Expected: {'Z': -1508}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000110; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 331,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1508
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100010; Y = 7'b1010010; // Expected: {'Z': -1564}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100010; Y = 7'b1010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 332,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1564
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b0110000; // Expected: {'Z': 2160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b0110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 333,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b1110100; // Expected: {'Z': 360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 334,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b1101010; // Expected: {'Z': 1386}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b1101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 335,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1386
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b0010111; // Expected: {'Z': 1196}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b0010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 336,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000011; Y = 7'b0100011; // Expected: {'Z': -2135}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000011; Y = 7'b0100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 337,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b1110000; // Expected: {'Z': 288}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 338,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011101; Y = 7'b0000010; // Expected: {'Z': -70}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011101; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 339,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101000; Y = 7'b1111001; // Expected: {'Z': -280}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101000; Y = 7'b1111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 340,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b1110111; // Expected: {'Z': -477}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b1110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 341,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -477
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111100; Y = 7'b1100100; // Expected: {'Z': -1680}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111100; Y = 7'b1100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 342,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010011; Y = 7'b1111100; // Expected: {'Z': 180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010011; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 343,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b1001101; // Expected: {'Z': 969}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b1001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 344,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 969
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001110; Y = 7'b1110100; // Expected: {'Z': 600}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001110; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 345,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b0100110; // Expected: {'Z': -1368}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 346,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b0001001; // Expected: {'Z': -306}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b0001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 347,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -306
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100011; Y = 7'b0110110; // Expected: {'Z': -1566}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100011; Y = 7'b0110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 348,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1566
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100011; Y = 7'b0010100; // Expected: {'Z': 700}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100011; Y = 7'b0010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 349,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101100; Y = 7'b0010111; // Expected: {'Z': 1012}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101100; Y = 7'b0010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 350,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1012
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000100; Y = 7'b1111110; // Expected: {'Z': 120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000100; Y = 7'b1111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 351,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110101; Y = 7'b0000010; // Expected: {'Z': -22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110101; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 352,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b0011011; // Expected: {'Z': -540}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b0011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 353,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011010; Y = 7'b0111010; // Expected: {'Z': -2204}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011010; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 354,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111001; Y = 7'b1100111; // Expected: {'Z': 175}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111001; Y = 7'b1100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 355,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b1010100; // Expected: {'Z': -880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b1010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 356,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011100; Y = 7'b1111101; // Expected: {'Z': -84}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011100; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 357,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b0111011; // Expected: {'Z': 1003}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 358,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1003
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000101; Y = 7'b1011011; // Expected: {'Z': -185}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000101; Y = 7'b1011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 359,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b0000101; // Expected: {'Z': 45}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b0000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 360,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100001; Y = 7'b0110000; // Expected: {'Z': 1584}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100001; Y = 7'b0110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 361,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1584
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011010; Y = 7'b0011011; // Expected: {'Z': 702}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011010; Y = 7'b0011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 362,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 702
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b0010011; // Expected: {'Z': 399}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b0010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 363,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 399
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101110; Y = 7'b0001101; // Expected: {'Z': 598}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101110; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 364,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 598
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111000; Y = 7'b1010111; // Expected: {'Z': -2296}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111000; Y = 7'b1010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 365,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000111; Y = 7'b1100001; // Expected: {'Z': 1767}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000111; Y = 7'b1100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 366,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1767
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b0011100; // Expected: {'Z': 476}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b0011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 367,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 476
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001011; Y = 7'b0110011; // Expected: {'Z': -2703}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001011; Y = 7'b0110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 368,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2703
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100101; Y = 7'b0111000; // Expected: {'Z': -1512}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100101; Y = 7'b0111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 369,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1512
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b1001110; // Expected: {'Z': 50}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b1001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 370,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111101; Y = 7'b0001101; // Expected: {'Z': 793}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111101; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 371,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 793
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b1010111; // Expected: {'Z': 2583}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b1010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 372,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2583
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110111; Y = 7'b1110011; // Expected: {'Z': -715}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110111; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 373,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -715
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000111; Y = 7'b0001000; // Expected: {'Z': -456}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000111; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 374,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001111; Y = 7'b0101101; // Expected: {'Z': -2205}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001111; Y = 7'b0101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 375,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101000; Y = 7'b1110101; // Expected: {'Z': 264}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101000; Y = 7'b1110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 376,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101000; Y = 7'b1101110; // Expected: {'Z': 432}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101000; Y = 7'b1101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 377,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110110; Y = 7'b1100101; // Expected: {'Z': -1458}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110110; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 378,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1458
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b1001001; // Expected: {'Z': -3410}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b1001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 379,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3410
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001001; Y = 7'b1101001; // Expected: {'Z': 1265}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001001; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 380,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1265
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001010; Y = 7'b0111001; // Expected: {'Z': 570}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001010; Y = 7'b0111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 381,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 570
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010001; Y = 7'b0011001; // Expected: {'Z': -1175}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010001; Y = 7'b0011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 382,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110000; Y = 7'b0100101; // Expected: {'Z': 1776}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110000; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 383,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1776
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b1011101; // Expected: {'Z': -1855}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b1011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 384,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1855
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101000; Y = 7'b0001101; // Expected: {'Z': -312}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101000; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 385,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -312
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100111; Y = 7'b1100001; // Expected: {'Z': 775}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100111; Y = 7'b1100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 386,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 775
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b0110011; // Expected: {'Z': -612}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b0110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 387,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010010; Y = 7'b0001111; // Expected: {'Z': -690}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010010; Y = 7'b0001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 388,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -690
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100000; Y = 7'b0000001; // Expected: {'Z': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100000; Y = 7'b0000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 389,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b1100110; // Expected: {'Z': 1248}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b1100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 390,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101110; Y = 7'b1011011; // Expected: {'Z': -1702}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101110; Y = 7'b1011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 391,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1702
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010011; Y = 7'b1110101; // Expected: {'Z': 495}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010011; Y = 7'b1110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 392,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 495
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100110; Y = 7'b0010110; // Expected: {'Z': 836}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100110; Y = 7'b0010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 393,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 836
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b0000101; // Expected: {'Z': 310}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b0000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 394,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 310
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000110; Y = 7'b1110011; // Expected: {'Z': -78}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000110; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 395,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110101; Y = 7'b1010111; // Expected: {'Z': 451}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110101; Y = 7'b1010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 396,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 451
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b1001011; // Expected: {'Z': 636}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b1001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 397,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 636
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101000; Y = 7'b1110011; // Expected: {'Z': -520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101000; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 398,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111101; Y = 7'b1010011; // Expected: {'Z': -2745}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111101; Y = 7'b1010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 399,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2745
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b1011011; // Expected: {'Z': 370}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b1011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 400,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 370
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010111; Y = 7'b0101100; // Expected: {'Z': 1012}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010111; Y = 7'b0101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 401,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1012
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101010; Y = 7'b0110100; // Expected: {'Z': 2184}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101010; Y = 7'b0110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 402,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b0010101; // Expected: {'Z': -714}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b0010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 403,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -714
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010011; Y = 7'b1110011; // Expected: {'Z': -247}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010011; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 404,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b1101110; // Expected: {'Z': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b1101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 405,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000111; Y = 7'b0010101; // Expected: {'Z': 147}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000111; Y = 7'b0010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 406,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b1111000; // Expected: {'Z': 96}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b1111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 407,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b0111011; // Expected: {'Z': -1888}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 408,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b0100010; // Expected: {'Z': 578}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b0100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 409,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 578
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111100; Y = 7'b0101111; // Expected: {'Z': -188}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111100; Y = 7'b0101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 410,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011010; Y = 7'b1011101; // Expected: {'Z': -910}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011010; Y = 7'b1011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 411,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -910
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b1101100; // Expected: {'Z': 1260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b1101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 412,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110001; Y = 7'b0000110; // Expected: {'Z': 294}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110001; Y = 7'b0000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 413,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 294
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b1010100; // Expected: {'Z': 748}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b1010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 414,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 748
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b0010010; // Expected: {'Z': -54}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b0010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 415,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001010; Y = 7'b1111000; // Expected: {'Z': 432}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001010; Y = 7'b1111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 416,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110000; Y = 7'b1011111; // Expected: {'Z': -1584}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110000; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 417,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1584
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000110; Y = 7'b1111101; // Expected: {'Z': -18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000110; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 418,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111000; Y = 7'b0001000; // Expected: {'Z': 448}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111000; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 419,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 448
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100101; Y = 7'b0000101; // Expected: {'Z': -135}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100101; Y = 7'b0000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 420,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010011; Y = 7'b0101111; // Expected: {'Z': -2115}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010011; Y = 7'b0101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 421,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2115
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001100; Y = 7'b1110000; // Expected: {'Z': 832}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001100; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 422,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 832
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001011; Y = 7'b0100000; // Expected: {'Z': -1696}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001011; Y = 7'b0100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 423,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1696
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001100; Y = 7'b0010110; // Expected: {'Z': -1144}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001100; Y = 7'b0010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 424,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111100; Y = 7'b0011010; // Expected: {'Z': 1560}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111100; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 425,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b0100110; // Expected: {'Z': -1216}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 426,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001000; Y = 7'b0000010; // Expected: {'Z': -112}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001000; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 427,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000111; Y = 7'b0000010; // Expected: {'Z': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000111; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 428,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b1011010; // Expected: {'Z': 1596}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b1011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 429,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1596
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000100; Y = 7'b1010110; // Expected: {'Z': -168}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000100; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 430,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110111; Y = 7'b1110001; // Expected: {'Z': -825}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110111; Y = 7'b1110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 431,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -825
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b0100101; // Expected: {'Z': -1036}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 432,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1036
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b1010101; // Expected: {'Z': -387}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b1010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 433,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -387
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100101; Y = 7'b0000011; // Expected: {'Z': 111}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100101; Y = 7'b0000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 434,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 111
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000011; Y = 7'b0000100; // Expected: {'Z': -244}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000011; Y = 7'b0000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 435,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b1000101; // Expected: {'Z': 1062}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b1000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 436,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1062
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110111; Y = 7'b1110000; // Expected: {'Z': 144}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110111; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 437,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b0101010; // Expected: {'Z': -1680}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b0101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 438,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b1110000; // Expected: {'Z': -16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 439,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001110; Y = 7'b0000111; // Expected: {'Z': -350}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001110; Y = 7'b0000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 440,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001110; Y = 7'b0111100; // Expected: {'Z': 840}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001110; Y = 7'b0111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 441,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110110; Y = 7'b1010011; // Expected: {'Z': -2430}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110110; Y = 7'b1010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 442,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b0110001; // Expected: {'Z': 833}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b0110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 443,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 833
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011111; Y = 7'b1011011; // Expected: {'Z': -1147}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011111; Y = 7'b1011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 444,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b1100010; // Expected: {'Z': -30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 445,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100101; Y = 7'b1010000; // Expected: {'Z': 1296}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100101; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 446,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b1111100; // Expected: {'Z': 76}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 447,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001101; Y = 7'b1001000; // Expected: {'Z': -728}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001101; Y = 7'b1001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 448,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100000; Y = 7'b0100110; // Expected: {'Z': 1216}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100000; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 449,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110110; Y = 7'b0010101; // Expected: {'Z': 1134}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110110; Y = 7'b0010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 450,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011010; Y = 7'b1101110; // Expected: {'Z': -468}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011010; Y = 7'b1101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 451,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -468
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001101; Y = 7'b1100010; // Expected: {'Z': -390}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001101; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 452,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -390
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b1010010; // Expected: {'Z': 1564}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b1010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 453,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1564
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101111; Y = 7'b0010000; // Expected: {'Z': 752}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101111; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 454,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 752
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b1001101; // Expected: {'Z': 612}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b1001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 455,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010010; Y = 7'b1110110; // Expected: {'Z': 460}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010010; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 456,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 460
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101111; Y = 7'b1000010; // Expected: {'Z': -2914}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101111; Y = 7'b1000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 457,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2914
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b0011101; // Expected: {'Z': 1305}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 458,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1305
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011010; Y = 7'b1110010; // Expected: {'Z': 532}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011010; Y = 7'b1110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 459,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 532
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000000; Y = 7'b0011010; // Expected: {'Z': -1664}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000000; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 460,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1664
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b0010100; // Expected: {'Z': 180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b0010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 461,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b1110000; // Expected: {'Z': 48}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 462,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000111; Y = 7'b0111100; // Expected: {'Z': -3420}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000111; Y = 7'b0111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 463,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001000; Y = 7'b1111110; // Expected: {'Z': -16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001000; Y = 7'b1111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 464,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011101; Y = 7'b0111111; // Expected: {'Z': -2205}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011101; Y = 7'b0111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 465,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100001; Y = 7'b1100010; // Expected: {'Z': 930}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100001; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 466,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 930
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111000; Y = 7'b0100011; // Expected: {'Z': -280}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111000; Y = 7'b0100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 467,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b1100101; // Expected: {'Z': -648}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 468,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111101; Y = 7'b1100000; // Expected: {'Z': -1952}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111101; Y = 7'b1100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 469,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1952
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b1101110; // Expected: {'Z': -306}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b1101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 470,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -306
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001011; Y = 7'b0001010; // Expected: {'Z': -530}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001011; Y = 7'b0001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 471,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -530
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000011; Y = 7'b0110110; // Expected: {'Z': -3294}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000011; Y = 7'b0110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 472,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3294
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010000; Y = 7'b0001100; // Expected: {'Z': 192}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010000; Y = 7'b0001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 473,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001111; Y = 7'b1000101; // Expected: {'Z': 2891}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001111; Y = 7'b1000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 474,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2891
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100110; Y = 7'b1011100; // Expected: {'Z': 936}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100110; Y = 7'b1011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 475,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 936
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b0011111; // Expected: {'Z': 1612}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b0011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 476,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b1000101; // Expected: {'Z': 1121}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b1000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 477,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010111; Y = 7'b1110001; // Expected: {'Z': -345}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010111; Y = 7'b1110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 478,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -345
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b1110100; // Expected: {'Z': 504}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 479,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100000; Y = 7'b0100101; // Expected: {'Z': 1184}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100000; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 480,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111101; Y = 7'b1101011; // Expected: {'Z': -1281}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111101; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 481,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1281
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b0100111; // Expected: {'Z': -39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b0100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 482,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000111; Y = 7'b1001010; // Expected: {'Z': -378}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000111; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 483,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -378
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000000; Y = 7'b1001000; // Expected: {'Z': 3584}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000000; Y = 7'b1001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 484,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3584
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111011; Y = 7'b1001010; // Expected: {'Z': 270}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111011; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 485,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 270
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b1001000; // Expected: {'Z': 1120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b1001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 486,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b1010000; // Expected: {'Z': -144}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 487,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000010; Y = 7'b1001110; // Expected: {'Z': -100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000010; Y = 7'b1001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 488,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000000; Y = 7'b0101110; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000000; Y = 7'b0101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 489,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110010; Y = 7'b1101001; // Expected: {'Z': -1150}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110010; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 490,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b1100011; // Expected: {'Z': 1044}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b1100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 491,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1044
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100000; Y = 7'b0000110; // Expected: {'Z': 192}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100000; Y = 7'b0000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 492,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b1100101; // Expected: {'Z': 810}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 493,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 810
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b1100001; // Expected: {'Z': 713}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b1100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 494,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 713
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101011; Y = 7'b0010001; // Expected: {'Z': -357}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101011; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 495,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -357
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111000; Y = 7'b0011010; // Expected: {'Z': 1456}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111000; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 496,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b0010111; // Expected: {'Z': 207}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b0010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 497,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 207
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000101; Y = 7'b1011011; // Expected: {'Z': -185}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000101; Y = 7'b1011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 498,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101110; Y = 7'b0111101; // Expected: {'Z': 2806}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101110; Y = 7'b0111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 499,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2806
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100101; Y = 7'b1100010; // Expected: {'Z': -1110}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100101; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 500,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111100; Y = 7'b1011101; // Expected: {'Z': 140}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111100; Y = 7'b1011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 501,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001011; Y = 7'b1101101; // Expected: {'Z': -209}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001011; Y = 7'b1101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 502,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b0010011; // Expected: {'Z': -57}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b0010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 503,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001110; Y = 7'b0000111; // Expected: {'Z': -350}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001110; Y = 7'b0000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 504,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b0110100; // Expected: {'Z': -988}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b0110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 505,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -988
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100111; Y = 7'b1101101; // Expected: {'Z': -741}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100111; Y = 7'b1101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 506,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -741
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b1010001; // Expected: {'Z': -2444}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 507,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2444
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011001; Y = 7'b0010000; // Expected: {'Z': 400}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011001; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 508,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010110; Y = 7'b0011110; // Expected: {'Z': 660}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010110; Y = 7'b0011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 509,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b0101010; // Expected: {'Z': 126}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b0101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 510,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001101; Y = 7'b1000100; // Expected: {'Z': 3060}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001101; Y = 7'b1000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 511,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001010; Y = 7'b0010110; // Expected: {'Z': 220}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001010; Y = 7'b0010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 512,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b0011001; // Expected: {'Z': -850}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b0011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 513,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -850
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101001; Y = 7'b0110011; // Expected: {'Z': 2091}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101001; Y = 7'b0110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 514,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2091
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000011; Y = 7'b0000111; // Expected: {'Z': -427}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000011; Y = 7'b0000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 515,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -427
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010111; Y = 7'b0111100; // Expected: {'Z': 1380}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010111; Y = 7'b0111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 516,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1380
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000010; Y = 7'b0101001; // Expected: {'Z': -2542}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000010; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 517,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2542
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001011; Y = 7'b0000100; // Expected: {'Z': -212}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001011; Y = 7'b0000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 518,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001010; Y = 7'b0010001; // Expected: {'Z': -918}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001010; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 519,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -918
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110111; Y = 7'b0100101; // Expected: {'Z': 2035}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110111; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 520,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2035
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b1010101; // Expected: {'Z': -2666}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b1010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 521,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2666
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b0011011; // Expected: {'Z': -1080}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b0011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 522,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010110; Y = 7'b0110001; // Expected: {'Z': 1078}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010110; Y = 7'b0110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 523,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1078
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110000; Y = 7'b1101000; // Expected: {'Z': 384}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110000; Y = 7'b1101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 524,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 384
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101011; Y = 7'b0100011; // Expected: {'Z': -735}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101011; Y = 7'b0100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 525,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -735
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b1110000; // Expected: {'Z': 576}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 526,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100100; Y = 7'b0110001; // Expected: {'Z': 1764}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100100; Y = 7'b0110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 527,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1764
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111100; Y = 7'b1001111; // Expected: {'Z': -2940}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111100; Y = 7'b1001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 528,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2940
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001101; Y = 7'b1100011; // Expected: {'Z': -377}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001101; Y = 7'b1100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 529,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -377
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010000; Y = 7'b0101100; // Expected: {'Z': 704}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010000; Y = 7'b0101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 530,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 704
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000000; Y = 7'b0110111; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000000; Y = 7'b0110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 531,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111011; Y = 7'b0001111; // Expected: {'Z': 885}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111011; Y = 7'b0001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 532,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 885
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100011; Y = 7'b0011011; // Expected: {'Z': 945}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100011; Y = 7'b0011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 533,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 945
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111011; Y = 7'b0111101; // Expected: {'Z': 3599}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111011; Y = 7'b0111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 534,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3599
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010110; Y = 7'b1011100; // Expected: {'Z': -792}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010110; Y = 7'b1011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 535,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b1110110; // Expected: {'Z': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 536,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b1010010; // Expected: {'Z': 782}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b1010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 537,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 782
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011101; Y = 7'b1001000; // Expected: {'Z': 1960}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011101; Y = 7'b1001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 538,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000100; Y = 7'b1110110; // Expected: {'Z': -40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000100; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 539,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000010; Y = 7'b1011101; // Expected: {'Z': 2170}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000010; Y = 7'b1011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 540,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100001; Y = 7'b0111011; // Expected: {'Z': -1829}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100001; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 541,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1829
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100011; Y = 7'b1010000; // Expected: {'Z': 1392}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100011; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 542,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111100; Y = 7'b1010110; // Expected: {'Z': 168}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111100; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 543,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111001; Y = 7'b1100001; // Expected: {'Z': 217}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111001; Y = 7'b1100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 544,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110011; Y = 7'b0110100; // Expected: {'Z': 2652}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110011; Y = 7'b0110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 545,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2652
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100001; Y = 7'b0010101; // Expected: {'Z': 693}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100001; Y = 7'b0010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 546,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 693
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011011; Y = 7'b1001100; // Expected: {'Z': -1404}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011011; Y = 7'b1001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 547,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1404
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011111; Y = 7'b1101101; // Expected: {'Z': -589}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011111; Y = 7'b1101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 548,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -589
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101100; Y = 7'b1000011; // Expected: {'Z': -2684}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101100; Y = 7'b1000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 549,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2684
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000100; Y = 7'b0110010; // Expected: {'Z': -3000}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000100; Y = 7'b0110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 550,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011010; Y = 7'b1001100; // Expected: {'Z': 1976}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011010; Y = 7'b1001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 551,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1976
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010111; Y = 7'b0011101; // Expected: {'Z': 667}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010111; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 552,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 667
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010110; Y = 7'b0111000; // Expected: {'Z': 1232}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010110; Y = 7'b0111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 553,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001011; Y = 7'b0110111; // Expected: {'Z': 605}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001011; Y = 7'b0110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 554,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 605
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001100; Y = 7'b1101111; // Expected: {'Z': -204}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001100; Y = 7'b1101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 555,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011011; Y = 7'b0110011; // Expected: {'Z': -1887}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011011; Y = 7'b0110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 556,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1887
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b1011110; // Expected: {'Z': 1632}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b1011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 557,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1632
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b1111000; // Expected: {'Z': -424}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b1111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 558,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -424
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001000; Y = 7'b0110111; // Expected: {'Z': -3080}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001000; Y = 7'b0110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 559,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b0110000; // Expected: {'Z': 2544}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b0110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 560,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2544
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001111; Y = 7'b0011000; // Expected: {'Z': -1176}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001111; Y = 7'b0011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 561,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b0110101; // Expected: {'Z': -3339}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 562,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3339
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b0110101; // Expected: {'Z': -954}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 563,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -954
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b1101110; // Expected: {'Z': 720}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b1101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 564,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b0111010; // Expected: {'Z': -580}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 565,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000010; Y = 7'b1111110; // Expected: {'Z': 124}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000010; Y = 7'b1111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 566,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101000; Y = 7'b1000011; // Expected: {'Z': 1464}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101000; Y = 7'b1000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 567,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001010; Y = 7'b0101010; // Expected: {'Z': 420}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001010; Y = 7'b0101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 568,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b0000001; // Expected: {'Z': -3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b0000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 569,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000100; Y = 7'b1000100; // Expected: {'Z': 3600}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000100; Y = 7'b1000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 570,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001100; Y = 7'b1010100; // Expected: {'Z': 2288}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001100; Y = 7'b1010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 571,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111100; Y = 7'b0111000; // Expected: {'Z': 3360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111100; Y = 7'b0111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 572,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011111; Y = 7'b1000011; // Expected: {'Z': 2013}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011111; Y = 7'b1000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 573,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2013
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b0010100; // Expected: {'Z': -720}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b0010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 574,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001001; Y = 7'b0011011; // Expected: {'Z': -1485}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001001; Y = 7'b0011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 575,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1485
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b0000101; // Expected: {'Z': -140}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b0000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 576,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111001; Y = 7'b1111001; // Expected: {'Z': 49}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111001; Y = 7'b1111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 577,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000000; Y = 7'b0111100; // Expected: {'Z': -3840}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000000; Y = 7'b0111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 578,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000000; Y = 7'b0000111; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000000; Y = 7'b0000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 579,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b1110010; // Expected: {'Z': -742}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b1110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 580,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -742
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001010; Y = 7'b1011100; // Expected: {'Z': 1944}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001010; Y = 7'b1011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 581,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011010; Y = 7'b0001000; // Expected: {'Z': 208}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011010; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 582,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001101; Y = 7'b0011110; // Expected: {'Z': -1530}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001101; Y = 7'b0011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 583,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1530
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010010; Y = 7'b0111110; // Expected: {'Z': 1116}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010010; Y = 7'b0111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 584,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101111; Y = 7'b1010010; // Expected: {'Z': -2162}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101111; Y = 7'b1010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 585,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b0101111; // Expected: {'Z': 47}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b0101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 586,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011010; Y = 7'b1001010; // Expected: {'Z': -1404}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011010; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 587,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1404
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011101; Y = 7'b0110111; // Expected: {'Z': 1595}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011101; Y = 7'b0110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 588,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1595
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110010; Y = 7'b1100001; // Expected: {'Z': -1550}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110010; Y = 7'b1100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 589,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010110; Y = 7'b1101000; // Expected: {'Z': -528}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010110; Y = 7'b1101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 590,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100111; Y = 7'b0100101; // Expected: {'Z': -925}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100111; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 591,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -925
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b1100111; // Expected: {'Z': 1050}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b1100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 592,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100001; Y = 7'b0101110; // Expected: {'Z': 1518}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100001; Y = 7'b0101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 593,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1518
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110011; Y = 7'b1000101; // Expected: {'Z': 767}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110011; Y = 7'b1000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 594,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 767
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011101; Y = 7'b1011101; // Expected: {'Z': -1015}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011101; Y = 7'b1011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 595,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1015
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b1101011; // Expected: {'Z': 63}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 596,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011110; Y = 7'b0110011; // Expected: {'Z': 1530}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011110; Y = 7'b0110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 597,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1530
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010100; Y = 7'b0001100; // Expected: {'Z': -528}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010100; Y = 7'b0001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 598,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b1111110; // Expected: {'Z': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b1111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 599,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b1010011; // Expected: {'Z': 1620}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b1010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 600,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b0110000; // Expected: {'Z': 1152}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b0110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 601,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011001; Y = 7'b0010000; // Expected: {'Z': -624}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011001; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 602,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000000; Y = 7'b1100111; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000000; Y = 7'b1100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 603,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010001; Y = 7'b0011011; // Expected: {'Z': -1269}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010001; Y = 7'b0011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 604,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1269
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001000; Y = 7'b0111101; // Expected: {'Z': 488}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001000; Y = 7'b0111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 605,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000111; Y = 7'b1100010; // Expected: {'Z': -210}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000111; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 606,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110010; Y = 7'b0001110; // Expected: {'Z': 700}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110010; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 607,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b0011111; // Expected: {'Z': -1953}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b0011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 608,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1953
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001110; Y = 7'b1100000; // Expected: {'Z': 1600}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001110; Y = 7'b1100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 609,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100000; Y = 7'b1111110; // Expected: {'Z': -64}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100000; Y = 7'b1111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 610,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111111; Y = 7'b1011110; // Expected: {'Z': -2142}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111111; Y = 7'b1011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 611,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000101; Y = 7'b1010001; // Expected: {'Z': -235}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000101; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 612,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -235
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111011; Y = 7'b1000000; // Expected: {'Z': -3776}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111011; Y = 7'b1000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 613,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3776
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001110; Y = 7'b1100010; // Expected: {'Z': 1500}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001110; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 614,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111011; Y = 7'b0001100; // Expected: {'Z': 708}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111011; Y = 7'b0001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 615,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 708
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b1011101; // Expected: {'Z': 665}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b1011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 616,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 665
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101010; Y = 7'b0001011; // Expected: {'Z': -242}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101010; Y = 7'b0001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 617,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101110; Y = 7'b0110000; // Expected: {'Z': 2208}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101110; Y = 7'b0110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 618,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001111; Y = 7'b0101111; // Expected: {'Z': -2303}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001111; Y = 7'b0101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 619,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2303
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b0010011; // Expected: {'Z': -912}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b0010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 620,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -912
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110010; Y = 7'b0001110; // Expected: {'Z': -196}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110010; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 621,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000111; Y = 7'b1100011; // Expected: {'Z': 1653}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000111; Y = 7'b1100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 622,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1653
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011011; Y = 7'b0011010; // Expected: {'Z': 702}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011011; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 623,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 702
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001110; Y = 7'b1100101; // Expected: {'Z': -378}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001110; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 624,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -378
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b0100110; // Expected: {'Z': -1064}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 625,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1064
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000101; Y = 7'b0101110; // Expected: {'Z': -2714}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000101; Y = 7'b0101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 626,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2714
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110001; Y = 7'b0010101; // Expected: {'Z': 1029}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110001; Y = 7'b0010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 627,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1029
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000011; Y = 7'b0011101; // Expected: {'Z': -1769}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000011; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 628,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1769
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111010; Y = 7'b1101100; // Expected: {'Z': -1160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111010; Y = 7'b1101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 629,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001011; Y = 7'b1011011; // Expected: {'Z': 1961}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001011; Y = 7'b1011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 630,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1961
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001000; Y = 7'b1011101; // Expected: {'Z': -280}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001000; Y = 7'b1011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 631,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b1100010; // Expected: {'Z': 1200}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 632,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b0100001; // Expected: {'Z': -1188}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b0100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 633,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b0000010; // Expected: {'Z': 124}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 634,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011010; Y = 7'b0011101; // Expected: {'Z': 754}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011010; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 635,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 754
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110101; Y = 7'b0111100; // Expected: {'Z': -660}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110101; Y = 7'b0111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 636,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010000; Y = 7'b1110010; // Expected: {'Z': -224}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010000; Y = 7'b1110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 637,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110011; Y = 7'b0010011; // Expected: {'Z': 969}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110011; Y = 7'b0010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 638,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 969
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b1111001; // Expected: {'Z': 238}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b1111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 639,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110011; Y = 7'b0111110; // Expected: {'Z': 3162}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110011; Y = 7'b0111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 640,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100110; Y = 7'b0010100; // Expected: {'Z': -520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100110; Y = 7'b0010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 641,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000010; Y = 7'b0001000; // Expected: {'Z': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000010; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 642,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b0111000; // Expected: {'Z': 3472}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b0111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 643,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3472
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b0010100; // Expected: {'Z': -340}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b0010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 644,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011010; Y = 7'b1011000; // Expected: {'Z': -1040}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011010; Y = 7'b1011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 645,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010111; Y = 7'b1010101; // Expected: {'Z': 1763}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010111; Y = 7'b1010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 646,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1763
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111001; Y = 7'b1100101; // Expected: {'Z': 189}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111001; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 647,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001100; Y = 7'b0010001; // Expected: {'Z': -884}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001100; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 648,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -884
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b0010101; // Expected: {'Z': -210}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b0010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 649,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001100; Y = 7'b0011001; // Expected: {'Z': 300}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001100; Y = 7'b0011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 650,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111010; Y = 7'b0101100; // Expected: {'Z': -264}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111010; Y = 7'b0101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 651,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b0101000; // Expected: {'Z': 960}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b0101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 652,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100001; Y = 7'b0011011; // Expected: {'Z': 891}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100001; Y = 7'b0011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 653,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 891
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000000; Y = 7'b1100011; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000000; Y = 7'b1100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 654,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b0100000; // Expected: {'Z': -96}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b0100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 655,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111100; Y = 7'b1111010; // Expected: {'Z': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111100; Y = 7'b1111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 656,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b0111011; // Expected: {'Z': -708}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 657,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -708
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011110; Y = 7'b1001111; // Expected: {'Z': -1470}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011110; Y = 7'b1001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 658,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1470
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001100; Y = 7'b1101111; // Expected: {'Z': -204}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001100; Y = 7'b1101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 659,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010110; Y = 7'b0110000; // Expected: {'Z': 1056}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010110; Y = 7'b0110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 660,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1056
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110110; Y = 7'b1110111; // Expected: {'Z': -486}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110110; Y = 7'b1110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 661,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -486
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000000; Y = 7'b0011100; // Expected: {'Z': -1792}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000000; Y = 7'b0011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 662,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001111; Y = 7'b1110111; // Expected: {'Z': 441}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001111; Y = 7'b1110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 663,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 441
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000111; Y = 7'b0010101; // Expected: {'Z': 147}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000111; Y = 7'b0010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 664,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000011; Y = 7'b1101011; // Expected: {'Z': 1281}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000011; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 665,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1281
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b1001101; // Expected: {'Z': 1530}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b1001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 666,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1530
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011111; Y = 7'b0011010; // Expected: {'Z': 806}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011111; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 667,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 806
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100001; Y = 7'b0111100; // Expected: {'Z': 1980}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100001; Y = 7'b0111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 668,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b1111101; // Expected: {'Z': 144}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 669,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b0011011; // Expected: {'Z': -486}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b0011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 670,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -486
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011001; Y = 7'b1110101; // Expected: {'Z': -275}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011001; Y = 7'b1110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 671,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -275
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b1010110; // Expected: {'Z': 420}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 672,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b1100110; // Expected: {'Z': -26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b1100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 673,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110011; Y = 7'b1100000; // Expected: {'Z': 416}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110011; Y = 7'b1100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 674,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000100; Y = 7'b1010101; // Expected: {'Z': 2580}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000100; Y = 7'b1010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 675,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100000; Y = 7'b0001101; // Expected: {'Z': 416}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100000; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 676,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b0011010; // Expected: {'Z': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 677,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b1110010; // Expected: {'Z': 420}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b1110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 678,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b0111001; // Expected: {'Z': 3534}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b0111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 679,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3534
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110011; Y = 7'b1101010; // Expected: {'Z': 286}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110011; Y = 7'b1101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 680,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 286
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111010; Y = 7'b0011101; // Expected: {'Z': 1682}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111010; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 681,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1682
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111001; Y = 7'b0100110; // Expected: {'Z': -266}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111001; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 682,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -266
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001010; Y = 7'b0011101; // Expected: {'Z': 290}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001010; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 683,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 290
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000010; Y = 7'b0101000; // Expected: {'Z': 80}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000010; Y = 7'b0101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 684,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010001; Y = 7'b1101001; // Expected: {'Z': 1081}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010001; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 685,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1081
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010100; Y = 7'b0011111; // Expected: {'Z': -1364}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010100; Y = 7'b0011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 686,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010010; Y = 7'b1110111; // Expected: {'Z': 414}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010010; Y = 7'b1110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 687,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 414
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011111; Y = 7'b1000001; // Expected: {'Z': 2079}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011111; Y = 7'b1000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 688,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2079
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111100; Y = 7'b0000011; // Expected: {'Z': 180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111100; Y = 7'b0000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 689,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b0001000; // Expected: {'Z': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 690,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111010; Y = 7'b1000010; // Expected: {'Z': -3596}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111010; Y = 7'b1000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 691,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3596
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101011; Y = 7'b0100011; // Expected: {'Z': 1505}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101011; Y = 7'b0100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 692,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1505
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011111; Y = 7'b0000100; // Expected: {'Z': 124}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011111; Y = 7'b0000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 693,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b1001100; // Expected: {'Z': 2184}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b1001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 694,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100001; Y = 7'b1111101; // Expected: {'Z': 93}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100001; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 695,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000101; Y = 7'b0110000; // Expected: {'Z': 240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000101; Y = 7'b0110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 696,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b0001011; // Expected: {'Z': -253}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b0001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 697,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001011; Y = 7'b1000101; // Expected: {'Z': -649}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001011; Y = 7'b1000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 698,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -649
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011001; Y = 7'b1001011; // Expected: {'Z': 2067}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011001; Y = 7'b1001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 699,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2067
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110011; Y = 7'b0110000; // Expected: {'Z': 2448}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110011; Y = 7'b0110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 700,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2448
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000110; Y = 7'b1110110; // Expected: {'Z': -60}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000110; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 701,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100111; Y = 7'b0001011; // Expected: {'Z': 429}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100111; Y = 7'b0001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 702,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 429
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010000; Y = 7'b0011100; // Expected: {'Z': 448}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010000; Y = 7'b0011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 703,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 448
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b1111110; // Expected: {'Z': -124}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b1111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 704,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001000; Y = 7'b0110110; // Expected: {'Z': -3024}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001000; Y = 7'b0110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 705,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111000; Y = 7'b1000100; // Expected: {'Z': -3360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111000; Y = 7'b1000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 706,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b1110111; // Expected: {'Z': 180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b1110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 707,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b0001000; // Expected: {'Z': 360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 708,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101110; Y = 7'b0100110; // Expected: {'Z': 1748}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101110; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 709,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1748
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011110; Y = 7'b1101010; // Expected: {'Z': -660}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011110; Y = 7'b1101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 710,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110111; Y = 7'b0101000; // Expected: {'Z': 2200}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110111; Y = 7'b0101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 711,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010010; Y = 7'b1000110; // Expected: {'Z': -1044}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010010; Y = 7'b1000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 712,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1044
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001010; Y = 7'b1010001; // Expected: {'Z': 2538}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001010; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 713,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2538
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000101; Y = 7'b1000001; // Expected: {'Z': 3717}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000101; Y = 7'b1000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 714,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3717
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001101; Y = 7'b0010000; // Expected: {'Z': -816}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001101; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 715,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b0001101; // Expected: {'Z': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 716,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011100; Y = 7'b1000110; // Expected: {'Z': -1624}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011100; Y = 7'b1000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 717,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b1101101; // Expected: {'Z': 285}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b1101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 718,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 285
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011010; Y = 7'b1011011; // Expected: {'Z': 1406}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011010; Y = 7'b1011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 719,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1406
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111111; Y = 7'b1011000; // Expected: {'Z': -2520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111111; Y = 7'b1011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 720,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b0000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b0000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 721,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b0000101; // Expected: {'Z': -315}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b0000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 722,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -315
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110000; Y = 7'b1011010; // Expected: {'Z': -1824}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110000; Y = 7'b1011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 723,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1824
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101010; Y = 7'b0100001; // Expected: {'Z': 1386}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101010; Y = 7'b0100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 724,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1386
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010011; Y = 7'b0001100; // Expected: {'Z': -540}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010011; Y = 7'b0001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 725,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000111; Y = 7'b1100000; // Expected: {'Z': 1824}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000111; Y = 7'b1100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 726,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1824
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111000; Y = 7'b1100001; // Expected: {'Z': 248}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111000; Y = 7'b1100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 727,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001011; Y = 7'b1011000; // Expected: {'Z': 2120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001011; Y = 7'b1011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 728,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011110; Y = 7'b1011111; // Expected: {'Z': -990}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011110; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 729,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -990
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010111; Y = 7'b0001011; // Expected: {'Z': 253}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010111; Y = 7'b0001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 730,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b1011011; // Expected: {'Z': 370}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b1011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 731,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 370
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000000; Y = 7'b1111101; // Expected: {'Z': 192}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000000; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 732,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011111; Y = 7'b0000010; // Expected: {'Z': -66}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011111; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 733,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000101; Y = 7'b0110000; // Expected: {'Z': -2832}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000101; Y = 7'b0110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 734,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2832
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000110; Y = 7'b1001001; // Expected: {'Z': -330}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000110; Y = 7'b1001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 735,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -330
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110010; Y = 7'b1110110; // Expected: {'Z': -500}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110010; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 736,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b0111110; // Expected: {'Z': -1426}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b0111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 737,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1426
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000100; Y = 7'b0110100; // Expected: {'Z': 208}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000100; Y = 7'b0110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 738,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000010; Y = 7'b0101011; // Expected: {'Z': 86}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000010; Y = 7'b0101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 739,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001110; Y = 7'b0100110; // Expected: {'Z': 532}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001110; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 740,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 532
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011011; Y = 7'b1100111; // Expected: {'Z': -675}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011011; Y = 7'b1100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 741,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -675
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b0001000; // Expected: {'Z': 424}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 742,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 424
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001111; Y = 7'b1111000; // Expected: {'Z': -120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001111; Y = 7'b1111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 743,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b1101000; // Expected: {'Z': 456}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b1101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 744,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011001; Y = 7'b0001001; // Expected: {'Z': -351}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011001; Y = 7'b0001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 745,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -351
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100010; Y = 7'b1001001; // Expected: {'Z': -1870}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100010; Y = 7'b1001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 746,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1870
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b0000111; // Expected: {'Z': 371}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b0000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 747,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 371
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b1101011; // Expected: {'Z': -420}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 748,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111010; Y = 7'b0110011; // Expected: {'Z': -306}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111010; Y = 7'b0110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 749,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -306
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000111; Y = 7'b0001101; // Expected: {'Z': -741}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000111; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 750,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -741
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b1101010; // Expected: {'Z': 506}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b1101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 751,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 506
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b0000010; // Expected: {'Z': -20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 752,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001000; Y = 7'b1111111; // Expected: {'Z': 56}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001000; Y = 7'b1111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 753,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110001; Y = 7'b0001000; // Expected: {'Z': 392}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110001; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 754,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b0011111; // Expected: {'Z': -1953}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b0011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 755,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1953
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011011; Y = 7'b0000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011011; Y = 7'b0000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 756,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b0000101; // Expected: {'Z': -95}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b0000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 757,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101011; Y = 7'b1111001; // Expected: {'Z': -301}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101011; Y = 7'b1111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 758,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -301
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b1111000; // Expected: {'Z': -360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b1111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 759,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001110; Y = 7'b1110000; // Expected: {'Z': -224}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001110; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 760,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001111; Y = 7'b0011100; // Expected: {'Z': 420}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001111; Y = 7'b0011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 761,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100110; Y = 7'b0011001; // Expected: {'Z': 950}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100110; Y = 7'b0011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 762,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b1010010; // Expected: {'Z': 1058}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b1010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 763,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1058
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100011; Y = 7'b1111110; // Expected: {'Z': 58}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100011; Y = 7'b1111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 764,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111110; Y = 7'b1010101; // Expected: {'Z': 86}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111110; Y = 7'b1010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 765,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b1101101; // Expected: {'Z': 646}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b1101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 766,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 646
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b1101100; // Expected: {'Z': -900}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b1101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 767,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011101; Y = 7'b1101011; // Expected: {'Z': -609}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011101; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 768,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -609
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001110; Y = 7'b0110100; // Expected: {'Z': -2600}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001110; Y = 7'b0110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 769,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011101; Y = 7'b1001100; // Expected: {'Z': 1820}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011101; Y = 7'b1001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 770,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110010; Y = 7'b1110011; // Expected: {'Z': -650}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110010; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 771,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b0100110; // Expected: {'Z': -38}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 772,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b1010110; // Expected: {'Z': 756}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 773,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011001; Y = 7'b0010010; // Expected: {'Z': -702}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011001; Y = 7'b0010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 774,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -702
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000010; Y = 7'b1001110; // Expected: {'Z': 3100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000010; Y = 7'b1001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 775,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001001; Y = 7'b0001110; // Expected: {'Z': -770}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001001; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 776,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -770
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000000; Y = 7'b0001110; // Expected: {'Z': -896}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000000; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 777,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b1000100; // Expected: {'Z': 600}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b1000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 778,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111010; Y = 7'b0100000; // Expected: {'Z': -192}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111010; Y = 7'b0100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 779,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b1001110; // Expected: {'Z': -150}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b1001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 780,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b0100011; // Expected: {'Z': -105}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b0100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 781,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001010; Y = 7'b0100110; // Expected: {'Z': -2052}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001010; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 782,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2052
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b0111011; // Expected: {'Z': -1003}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 783,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1003
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b1001111; // Expected: {'Z': 3087}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b1001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 784,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3087
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101011; Y = 7'b1000010; // Expected: {'Z': -2666}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101011; Y = 7'b1000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 785,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2666
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110001; Y = 7'b1110000; // Expected: {'Z': -784}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110001; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 786,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011010; Y = 7'b1011111; // Expected: {'Z': -858}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011010; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 787,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -858
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000101; Y = 7'b0111000; // Expected: {'Z': -3304}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000101; Y = 7'b0111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 788,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3304
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001010; Y = 7'b0101011; // Expected: {'Z': 430}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001010; Y = 7'b0101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 789,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110010; Y = 7'b0011101; // Expected: {'Z': 1450}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110010; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 790,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001110; Y = 7'b1000100; // Expected: {'Z': -840}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001110; Y = 7'b1000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 791,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b1011010; // Expected: {'Z': -114}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b1011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 792,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000010; Y = 7'b1000110; // Expected: {'Z': -116}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000010; Y = 7'b1000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 793,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110001; Y = 7'b1111011; // Expected: {'Z': -245}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110001; Y = 7'b1111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 794,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000000; Y = 7'b1011010; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000000; Y = 7'b1011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 795,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110111; Y = 7'b0100011; // Expected: {'Z': 1925}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110111; Y = 7'b0100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 796,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1925
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110000; Y = 7'b0001111; // Expected: {'Z': -240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110000; Y = 7'b0001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 797,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b0101110; // Expected: {'Z': -874}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b0101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 798,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -874
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101111; Y = 7'b0000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101111; Y = 7'b0000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 799,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b1101000; // Expected: {'Z': 960}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b1101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 800,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010111; Y = 7'b1001011; // Expected: {'Z': -1219}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010111; Y = 7'b1001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 801,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1219
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b0111111; // Expected: {'Z': -1890}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b0111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 802,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1890
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111011; Y = 7'b1110000; // Expected: {'Z': 80}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111011; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 803,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101011; Y = 7'b1001111; // Expected: {'Z': -2107}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101011; Y = 7'b1001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 804,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b1010110; // Expected: {'Z': 2646}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 805,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2646
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b1010001; // Expected: {'Z': 141}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 806,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011011; Y = 7'b1111111; // Expected: {'Z': 37}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011011; Y = 7'b1111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 807,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110001; Y = 7'b1110100; // Expected: {'Z': -588}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110001; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 808,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -588
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001001; Y = 7'b1000010; // Expected: {'Z': 3410}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001001; Y = 7'b1000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 809,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3410
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101011; Y = 7'b0011011; // Expected: {'Z': -567}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101011; Y = 7'b0011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 810,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -567
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001100; Y = 7'b1011100; // Expected: {'Z': -432}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001100; Y = 7'b1011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 811,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010111; Y = 7'b1000100; // Expected: {'Z': -1380}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010111; Y = 7'b1000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 812,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1380
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100110; Y = 7'b1100011; // Expected: {'Z': -1102}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100110; Y = 7'b1100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 813,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b0101110; // Expected: {'Z': -1472}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b0101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 814,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1472
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b0011001; // Expected: {'Z': -450}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b0011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 815,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010111; Y = 7'b1001000; // Expected: {'Z': 2296}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010111; Y = 7'b1001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 816,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110011; Y = 7'b0100111; // Expected: {'Z': 1989}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110011; Y = 7'b0100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 817,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1989
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b0000010; // Expected: {'Z': -6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 818,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111100; Y = 7'b0011010; // Expected: {'Z': 1560}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111100; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 819,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b0101011; // Expected: {'Z': -1204}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b0101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 820,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100111; Y = 7'b1011101; // Expected: {'Z': 875}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100111; Y = 7'b1011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 821,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 875
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b1010100; // Expected: {'Z': 1584}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b1010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 822,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1584
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011100; Y = 7'b1011010; // Expected: {'Z': -1064}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011100; Y = 7'b1011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 823,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1064
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101010; Y = 7'b1110110; // Expected: {'Z': -420}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101010; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 824,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b0001000; // Expected: {'Z': -288}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 825,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000111; Y = 7'b1001111; // Expected: {'Z': -343}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000111; Y = 7'b1001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 826,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -343
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010010; Y = 7'b0010000; // Expected: {'Z': -736}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010010; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 827,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101000; Y = 7'b0010010; // Expected: {'Z': 720}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101000; Y = 7'b0010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 828,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001011; Y = 7'b0011100; // Expected: {'Z': -1484}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001011; Y = 7'b0011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 829,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1484
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010111; Y = 7'b1100001; // Expected: {'Z': 1271}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010111; Y = 7'b1100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 830,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1271
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111101; Y = 7'b1001110; // Expected: {'Z': -3050}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111101; Y = 7'b1001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 831,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111010; Y = 7'b1001111; // Expected: {'Z': 294}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111010; Y = 7'b1001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 832,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 294
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101010; Y = 7'b0101011; // Expected: {'Z': -946}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101010; Y = 7'b0101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 833,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -946
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b0010111; // Expected: {'Z': 1426}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b0010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 834,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1426
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b0000001; // Expected: {'Z': -23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b0000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 835,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100000; Y = 7'b1000100; // Expected: {'Z': -1920}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100000; Y = 7'b1000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 836,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b1100011; // Expected: {'Z': 580}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b1100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 837,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b1011110; // Expected: {'Z': -680}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b1011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 838,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010011; Y = 7'b1111010; // Expected: {'Z': 270}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010011; Y = 7'b1111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 839,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 270
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110111; Y = 7'b0101000; // Expected: {'Z': -360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110111; Y = 7'b0101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 840,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b0010101; // Expected: {'Z': -672}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b0010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 841,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100011; Y = 7'b0010011; // Expected: {'Z': 665}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100011; Y = 7'b0010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 842,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 665
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b1001000; // Expected: {'Z': -1176}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b1001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 843,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111101; Y = 7'b0111100; // Expected: {'Z': 3660}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111101; Y = 7'b0111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 844,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b1101010; // Expected: {'Z': 704}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b1101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 845,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 704
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011011; Y = 7'b0100010; // Expected: {'Z': 918}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011011; Y = 7'b0100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 846,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 918
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010001; Y = 7'b1101000; // Expected: {'Z': 1128}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010001; Y = 7'b1101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 847,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110011; Y = 7'b0010001; // Expected: {'Z': 867}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110011; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 848,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 867
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110011; Y = 7'b1001010; // Expected: {'Z': 702}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110011; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 849,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 702
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001101; Y = 7'b1100000; // Expected: {'Z': 1632}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001101; Y = 7'b1100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 850,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1632
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b0001001; // Expected: {'Z': -162}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b0001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 851,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000100; Y = 7'b1101100; // Expected: {'Z': 1200}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000100; Y = 7'b1101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 852,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100001; Y = 7'b0001101; // Expected: {'Z': 429}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100001; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 853,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 429
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111111; Y = 7'b1111110; // Expected: {'Z': -126}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111111; Y = 7'b1111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 854,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b0001101; // Expected: {'Z': -364}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 855,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001000; Y = 7'b1100111; // Expected: {'Z': 1400}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001000; Y = 7'b1100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 856,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111111; Y = 7'b0111101; // Expected: {'Z': 3843}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111111; Y = 7'b0111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 857,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3843
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010111; Y = 7'b1000001; // Expected: {'Z': 2583}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010111; Y = 7'b1000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 858,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2583
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b0001110; // Expected: {'Z': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 859,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010001; Y = 7'b1101011; // Expected: {'Z': 987}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010001; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 860,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 987
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010010; Y = 7'b1010011; // Expected: {'Z': -810}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010010; Y = 7'b1010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 861,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -810
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b0101101; // Expected: {'Z': -855}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b0101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 862,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -855
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011100; Y = 7'b0100001; // Expected: {'Z': 924}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011100; Y = 7'b0100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 863,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 924
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100011; Y = 7'b0101110; // Expected: {'Z': 1610}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100011; Y = 7'b0101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 864,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1610
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b1010011; // Expected: {'Z': 765}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b1010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 865,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 765
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b0000001; // Expected: {'Z': -19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b0000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 866,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b0110001; // Expected: {'Z': 3038}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b0110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 867,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3038
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110111; Y = 7'b1110011; // Expected: {'Z': -715}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110111; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 868,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -715
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100101; Y = 7'b0111001; // Expected: {'Z': 2109}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100101; Y = 7'b0111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 869,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2109
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101100; Y = 7'b0101000; // Expected: {'Z': 1760}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101100; Y = 7'b0101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 870,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111101; Y = 7'b1100111; // Expected: {'Z': -1525}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111101; Y = 7'b1100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 871,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1525
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000111; Y = 7'b1111001; // Expected: {'Z': 399}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000111; Y = 7'b1111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 872,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 399
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001110; Y = 7'b1010001; // Expected: {'Z': 2350}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001110; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 873,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b0110110; // Expected: {'Z': -918}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b0110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 874,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -918
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011111; Y = 7'b0101101; // Expected: {'Z': -1485}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011111; Y = 7'b0101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 875,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1485
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b0001101; // Expected: {'Z': -364}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 876,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b0100001; // Expected: {'Z': -1122}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b0100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 877,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b0010111; // Expected: {'Z': 207}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b0010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 878,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 207
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b0110101; // Expected: {'Z': 901}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 879,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 901
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b1001101; // Expected: {'Z': 969}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b1001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 880,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 969
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010111; Y = 7'b1000001; // Expected: {'Z': -1449}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010111; Y = 7'b1000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 881,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1449
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100001; Y = 7'b1000101; // Expected: {'Z': -1947}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100001; Y = 7'b1000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 882,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1947
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111010; Y = 7'b0001100; // Expected: {'Z': 696}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111010; Y = 7'b0001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 883,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 696
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010111; Y = 7'b0100010; // Expected: {'Z': -1394}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010111; Y = 7'b0100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 884,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1394
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b0010000; // Expected: {'Z': 720}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 885,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100111; Y = 7'b0101011; // Expected: {'Z': -1075}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100111; Y = 7'b0101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 886,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1075
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000010; Y = 7'b1000111; // Expected: {'Z': 3534}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000010; Y = 7'b1000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 887,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3534
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010101; Y = 7'b0101101; // Expected: {'Z': -1935}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010101; Y = 7'b0101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 888,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1935
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b1100001; // Expected: {'Z': -527}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b1100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 889,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -527
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b0000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b0000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 890,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b1110011; // Expected: {'Z': 299}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 891,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 299
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011010; Y = 7'b0010010; // Expected: {'Z': -684}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011010; Y = 7'b0010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 892,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -684
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b0001001; // Expected: {'Z': -324}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b0001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 893,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -324
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b1000001; // Expected: {'Z': 630}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b1000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 894,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 630
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b1000011; // Expected: {'Z': 2440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b1000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 895,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100101; Y = 7'b0100100; // Expected: {'Z': -972}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100101; Y = 7'b0100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 896,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -972
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100110; Y = 7'b0001100; // Expected: {'Z': -312}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100110; Y = 7'b0001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 897,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -312
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101011; Y = 7'b1110110; // Expected: {'Z': 210}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101011; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 898,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000000; Y = 7'b1101100; // Expected: {'Z': 1280}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000000; Y = 7'b1101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 899,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001001; Y = 7'b0010110; // Expected: {'Z': -1210}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001001; Y = 7'b0010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 900,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101100; Y = 7'b0001000; // Expected: {'Z': 352}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101100; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 901,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001110; Y = 7'b1110001; // Expected: {'Z': 750}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001110; Y = 7'b1110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 902,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b1101001; // Expected: {'Z': 414}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 903,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 414
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110011; Y = 7'b1110110; // Expected: {'Z': 130}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110011; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 904,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100111; Y = 7'b0101000; // Expected: {'Z': 1560}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100111; Y = 7'b0101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 905,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110011; Y = 7'b1010001; // Expected: {'Z': 611}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110011; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 906,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 611
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010101; Y = 7'b1010101; // Expected: {'Z': 1849}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010101; Y = 7'b1010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 907,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1849
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b0111101; // Expected: {'Z': -1037}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b0111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 908,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1037
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100111; Y = 7'b0101111; // Expected: {'Z': -1175}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100111; Y = 7'b0101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 909,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111011; Y = 7'b0000100; // Expected: {'Z': -20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111011; Y = 7'b0000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 910,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b1010011; // Expected: {'Z': 540}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b1010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 911,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001000; Y = 7'b0101100; // Expected: {'Z': 352}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001000; Y = 7'b0101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 912,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000000; Y = 7'b0000010; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000000; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 913,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b1001010; // Expected: {'Z': 2268}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 914,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2268
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001111; Y = 7'b1010111; // Expected: {'Z': 2009}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001111; Y = 7'b1010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 915,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2009
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001010; Y = 7'b1011100; // Expected: {'Z': -360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001010; Y = 7'b1011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 916,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111010; Y = 7'b0001001; // Expected: {'Z': -54}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111010; Y = 7'b0001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 917,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010011; Y = 7'b1001110; // Expected: {'Z': 2250}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010011; Y = 7'b1001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 918,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b0000101; // Expected: {'Z': -200}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b0000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 919,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b1110011; // Expected: {'Z': 156}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 920,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011001; Y = 7'b0110100; // Expected: {'Z': -2028}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011001; Y = 7'b0110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 921,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2028
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010000; Y = 7'b0001000; // Expected: {'Z': 128}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010000; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 922,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b0001011; // Expected: {'Z': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b0001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 923,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b1100101; // Expected: {'Z': 621}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 924,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 621
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001000; Y = 7'b0111100; // Expected: {'Z': -3360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001000; Y = 7'b0111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 925,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101011; Y = 7'b1000101; // Expected: {'Z': -2537}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101011; Y = 7'b1000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 926,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2537
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110001; Y = 7'b0001000; // Expected: {'Z': 392}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110001; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 927,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b1110000; // Expected: {'Z': 544}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 928,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 544
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000011; Y = 7'b0000101; // Expected: {'Z': -305}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000011; Y = 7'b0000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 929,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -305
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011011; Y = 7'b1111111; // Expected: {'Z': -27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011011; Y = 7'b1111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 930,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111010; Y = 7'b0011100; // Expected: {'Z': 1624}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111010; Y = 7'b0011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 931,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110000; Y = 7'b1001001; // Expected: {'Z': 880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110000; Y = 7'b1001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 932,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100100; Y = 7'b0110101; // Expected: {'Z': 1908}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100100; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 933,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1908
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101011; Y = 7'b1101010; // Expected: {'Z': 462}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101011; Y = 7'b1101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 934,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000100; Y = 7'b1101111; // Expected: {'Z': 1020}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000100; Y = 7'b1101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 935,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1020
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b1011010; // Expected: {'Z': -2356}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b1011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 936,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2356
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101000; Y = 7'b1010000; // Expected: {'Z': -1920}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101000; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 937,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100111; Y = 7'b0100101; // Expected: {'Z': -925}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100111; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 938,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -925
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b0010110; // Expected: {'Z': -1386}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b0010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 939,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1386
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011011; Y = 7'b0010101; // Expected: {'Z': 567}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011011; Y = 7'b0010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 940,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 567
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001100; Y = 7'b0010000; // Expected: {'Z': -832}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001100; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 941,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -832
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b0010010; // Expected: {'Z': -756}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b0010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 942,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000100; Y = 7'b0111101; // Expected: {'Z': -3660}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000100; Y = 7'b0111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 943,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101001; Y = 7'b0111101; // Expected: {'Z': 2501}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101001; Y = 7'b0111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 944,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2501
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110111; Y = 7'b0000111; // Expected: {'Z': -63}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110111; Y = 7'b0000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 945,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b0110111; // Expected: {'Z': -1980}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b0110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 946,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001000; Y = 7'b0010100; // Expected: {'Z': -1120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001000; Y = 7'b0010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 947,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b0011111; // Expected: {'Z': 620}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b0011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 948,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b0000001; // Expected: {'Z': -18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b0000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 949,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b1011000; // Expected: {'Z': 400}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b1011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 950,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b1100001; // Expected: {'Z': 372}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b1100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 951,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 372
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100110; Y = 7'b1101010; // Expected: {'Z': 572}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100110; Y = 7'b1101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 952,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 572
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010011; Y = 7'b1110110; // Expected: {'Z': 450}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010011; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 953,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011111; Y = 7'b1100101; // Expected: {'Z': 891}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011111; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 954,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 891
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011001; Y = 7'b1001000; // Expected: {'Z': -1400}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011001; Y = 7'b1001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 955,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001100; Y = 7'b1101000; // Expected: {'Z': 1248}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001100; Y = 7'b1101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 956,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111000; Y = 7'b1101011; // Expected: {'Z': 168}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111000; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 957,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010011; Y = 7'b0111101; // Expected: {'Z': -2745}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010011; Y = 7'b0111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 958,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2745
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011111; Y = 7'b1000011; // Expected: {'Z': -1891}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011111; Y = 7'b1000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 959,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1891
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000011; Y = 7'b0010001; // Expected: {'Z': -1037}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000011; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 960,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1037
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b0101001; // Expected: {'Z': -779}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 961,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -779
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111100; Y = 7'b0000010; // Expected: {'Z': 120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111100; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 962,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011110; Y = 7'b1100111; // Expected: {'Z': -750}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011110; Y = 7'b1100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 963,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011110; Y = 7'b0110101; // Expected: {'Z': 1590}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011110; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 964,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1590
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010100; Y = 7'b0100001; // Expected: {'Z': -1452}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010100; Y = 7'b0100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 965,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1452
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b1001000; // Expected: {'Z': 1680}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b1001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 966,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010100; Y = 7'b1110101; // Expected: {'Z': 484}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010100; Y = 7'b1110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 967,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 484
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010011; Y = 7'b0100100; // Expected: {'Z': 684}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010011; Y = 7'b0100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 968,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 684
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000111; Y = 7'b0001111; // Expected: {'Z': -855}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000111; Y = 7'b0001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 969,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -855
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011001; Y = 7'b0010000; // Expected: {'Z': 400}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011001; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 970,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110010; Y = 7'b0100110; // Expected: {'Z': -532}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110010; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 971,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -532
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111110; Y = 7'b0111001; // Expected: {'Z': -114}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111110; Y = 7'b0111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 972,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100101; Y = 7'b1110011; // Expected: {'Z': -481}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100101; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 973,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -481
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111100; Y = 7'b1011111; // Expected: {'Z': -1980}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111100; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 974,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011001; Y = 7'b1010000; // Expected: {'Z': 1872}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011001; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 975,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1872
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111100; Y = 7'b0010101; // Expected: {'Z': -84}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111100; Y = 7'b0010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 976,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001110; Y = 7'b0111111; // Expected: {'Z': 882}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001110; Y = 7'b0111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 977,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 882
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011100; Y = 7'b1111000; // Expected: {'Z': -224}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011100; Y = 7'b1111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 978,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011100; Y = 7'b1001111; // Expected: {'Z': -1372}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011100; Y = 7'b1001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 979,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1372
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111100; Y = 7'b0011100; // Expected: {'Z': -112}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111100; Y = 7'b0011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 980,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000100; Y = 7'b1010101; // Expected: {'Z': -172}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000100; Y = 7'b1010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 981,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b1001100; // Expected: {'Z': 1664}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b1001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 982,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1664
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b0000001; // Expected: {'Z': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b0000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 983,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000010; Y = 7'b0011100; // Expected: {'Z': -1736}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000010; Y = 7'b0011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 984,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101011; Y = 7'b0110100; // Expected: {'Z': 2236}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101011; Y = 7'b0110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 985,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b0101001; // Expected: {'Z': -820}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 986,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b0011001; // Expected: {'Z': -575}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b0011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 987,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -575
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000110; Y = 7'b0110001; // Expected: {'Z': 294}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000110; Y = 7'b0110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 988,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 294
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111101; Y = 7'b1110100; // Expected: {'Z': -732}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111101; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 989,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -732
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110000; Y = 7'b0111101; // Expected: {'Z': -976}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110000; Y = 7'b0111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 990,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -976
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000111; Y = 7'b0101110; // Expected: {'Z': -2622}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000111; Y = 7'b0101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 991,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2622
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010000; Y = 7'b1110010; // Expected: {'Z': -224}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010000; Y = 7'b1110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 992,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001011; Y = 7'b1010100; // Expected: {'Z': -484}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001011; Y = 7'b1010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 993,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -484
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b1011101; // Expected: {'Z': -35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b1011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 994,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b0010001; // Expected: {'Z': 408}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 995,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001010; Y = 7'b1010010; // Expected: {'Z': -460}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001010; Y = 7'b1010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 996,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -460
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000111; Y = 7'b1101101; // Expected: {'Z': -133}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000111; Y = 7'b1101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 997,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -133
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111000; Y = 7'b0110110; // Expected: {'Z': 3024}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111000; Y = 7'b0110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 998,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110000; Y = 7'b1000011; // Expected: {'Z': -2928}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110000; Y = 7'b1000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 999,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2928
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b1111000; // Expected: {'Z': -496}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b1111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1000,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b0111010; // Expected: {'Z': -2784}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1001,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b0100100; // Expected: {'Z': -648}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b0100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1002,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b1011001; // Expected: {'Z': 1170}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b1011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1003,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010011; Y = 7'b0100001; // Expected: {'Z': -1485}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010011; Y = 7'b0100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1004,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1485
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011010; Y = 7'b1100010; // Expected: {'Z': 1140}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011010; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1005,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001010; Y = 7'b0001011; // Expected: {'Z': 110}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001010; Y = 7'b0001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1006,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111000; Y = 7'b0111010; // Expected: {'Z': -464}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111000; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1007,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110111; Y = 7'b0110011; // Expected: {'Z': -459}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110111; Y = 7'b0110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1008,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -459
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011011; Y = 7'b0010010; // Expected: {'Z': 486}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011011; Y = 7'b0010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1009,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 486
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111010; Y = 7'b0001101; // Expected: {'Z': 754}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111010; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1010,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 754
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010110; Y = 7'b1001110; // Expected: {'Z': -1100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010110; Y = 7'b1001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1011,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011011; Y = 7'b0111010; // Expected: {'Z': 1566}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011011; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1012,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1566
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111111; Y = 7'b1101011; // Expected: {'Z': -1323}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111111; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1013,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1323
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b0011000; // Expected: {'Z': -360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b0011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1014,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b1101111; // Expected: {'Z': 204}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b1101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1015,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001111; Y = 7'b0011001; // Expected: {'Z': 375}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001111; Y = 7'b0011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1016,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 375
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b0000111; // Expected: {'Z': -441}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b0000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1017,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -441
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010011; Y = 7'b0100011; // Expected: {'Z': -1575}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010011; Y = 7'b0100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1018,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1575
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b1010011; // Expected: {'Z': 1260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b1010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1019,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100100; Y = 7'b0010001; // Expected: {'Z': 612}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100100; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1020,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001011; Y = 7'b1100110; // Expected: {'Z': -286}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001011; Y = 7'b1100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1021,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -286
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111010; Y = 7'b0001111; // Expected: {'Z': -90}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111010; Y = 7'b0001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1022,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010010; Y = 7'b1100010; // Expected: {'Z': -540}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010010; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1023,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011011; Y = 7'b1101001; // Expected: {'Z': 851}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011011; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1024,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 851
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000110; Y = 7'b1011100; // Expected: {'Z': -216}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000110; Y = 7'b1011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1025,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010000; Y = 7'b0001010; // Expected: {'Z': 160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010000; Y = 7'b0001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1026,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010110; Y = 7'b0100011; // Expected: {'Z': 770}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010110; Y = 7'b0100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1027,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 770
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110001; Y = 7'b0001110; // Expected: {'Z': 686}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110001; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1028,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 686
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b0101101; // Expected: {'Z': -765}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b0101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1029,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -765
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011011; Y = 7'b1111011; // Expected: {'Z': 185}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011011; Y = 7'b1111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1030,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111100; Y = 7'b0010101; // Expected: {'Z': -84}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111100; Y = 7'b0010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1031,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111001; Y = 7'b1100111; // Expected: {'Z': 175}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111001; Y = 7'b1100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1032,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b1110100; // Expected: {'Z': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1033,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b0010011; // Expected: {'Z': -380}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b0010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1034,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -380
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111000; Y = 7'b1110000; // Expected: {'Z': 128}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111000; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1035,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100011; Y = 7'b0010101; // Expected: {'Z': 735}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100011; Y = 7'b0010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1036,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 735
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b1110010; // Expected: {'Z': 588}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b1110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1037,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 588
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001110; Y = 7'b0010000; // Expected: {'Z': 224}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001110; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1038,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100111; Y = 7'b0000100; // Expected: {'Z': 156}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100111; Y = 7'b0000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1039,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101111; Y = 7'b0110111; // Expected: {'Z': 2585}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101111; Y = 7'b0110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1040,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2585
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010010; Y = 7'b0100000; // Expected: {'Z': -1472}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010010; Y = 7'b0100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1041,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1472
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101010; Y = 7'b1000010; // Expected: {'Z': 1364}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101010; Y = 7'b1000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1042,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101011; Y = 7'b0001011; // Expected: {'Z': -231}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101011; Y = 7'b0001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1043,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111101; Y = 7'b0001110; // Expected: {'Z': 854}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111101; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1044,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 854
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000010; Y = 7'b1111111; // Expected: {'Z': -2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000010; Y = 7'b1111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1045,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000111; Y = 7'b0111011; // Expected: {'Z': 413}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000111; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1046,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 413
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100101; Y = 7'b1111010; // Expected: {'Z': -222}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100101; Y = 7'b1111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1047,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110110; Y = 7'b0000110; // Expected: {'Z': 324}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110110; Y = 7'b0000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1048,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 324
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000111; Y = 7'b0110100; // Expected: {'Z': 364}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000111; Y = 7'b0110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1049,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110000; Y = 7'b1011100; // Expected: {'Z': -1728}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110000; Y = 7'b1011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1050,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101000; Y = 7'b1110010; // Expected: {'Z': -560}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101000; Y = 7'b1110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1051,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000110; Y = 7'b1111101; // Expected: {'Z': 174}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000110; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1052,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001011; Y = 7'b1100100; // Expected: {'Z': 1484}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001011; Y = 7'b1100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1053,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1484
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110010; Y = 7'b1001110; // Expected: {'Z': 700}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110010; Y = 7'b1001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1054,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100111; Y = 7'b0110111; // Expected: {'Z': -1375}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100111; Y = 7'b0110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1055,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1375
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b1011100; // Expected: {'Z': 1008}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b1011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1056,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111011; Y = 7'b1110110; // Expected: {'Z': -590}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111011; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1057,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -590
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110111; Y = 7'b0010010; // Expected: {'Z': 990}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110111; Y = 7'b0010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1058,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 990
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010111; Y = 7'b0000010; // Expected: {'Z': -82}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010111; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1059,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -82
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011010; Y = 7'b0101101; // Expected: {'Z': -1710}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011010; Y = 7'b0101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1060,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1710
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000010; Y = 7'b1101011; // Expected: {'Z': 1302}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000010; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1061,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1302
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000110; Y = 7'b1000111; // Expected: {'Z': -342}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000110; Y = 7'b1000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1062,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -342
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101010; Y = 7'b1001111; // Expected: {'Z': 1078}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101010; Y = 7'b1001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1063,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1078
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100001; Y = 7'b0110101; // Expected: {'Z': -1643}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100001; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1064,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1643
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b0011111; // Expected: {'Z': -1054}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b0011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1065,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1054
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111000; Y = 7'b1100100; // Expected: {'Z': -1568}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111000; Y = 7'b1100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1066,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1568
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000110; Y = 7'b0001001; // Expected: {'Z': -522}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000110; Y = 7'b0001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1067,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -522
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b0011010; // Expected: {'Z': 1612}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1068,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100011; Y = 7'b0111001; // Expected: {'Z': -1653}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100011; Y = 7'b0111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1069,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1653
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b1110100; // Expected: {'Z': -108}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1070,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b0000011; // Expected: {'Z': -189}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b0000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1071,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b0001011; // Expected: {'Z': 495}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b0001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1072,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 495
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001100; Y = 7'b1000101; // Expected: {'Z': -708}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001100; Y = 7'b1000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1073,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -708
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111011; Y = 7'b1001100; // Expected: {'Z': 260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111011; Y = 7'b1001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1074,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b1110000; // Expected: {'Z': 48}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1075,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110111; Y = 7'b0101001; // Expected: {'Z': -369}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110111; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1076,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -369
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b0111011; // Expected: {'Z': 1180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1077,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b1111101; // Expected: {'Z': -186}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1078,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110111; Y = 7'b0100001; // Expected: {'Z': 1815}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110111; Y = 7'b0100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1079,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1815
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010010; Y = 7'b0010011; // Expected: {'Z': -874}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010010; Y = 7'b0010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1080,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -874
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001111; Y = 7'b1000001; // Expected: {'Z': -945}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001111; Y = 7'b1000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1081,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -945
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b1010111; // Expected: {'Z': -984}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b1010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1082,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -984
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111010; Y = 7'b1111000; // Expected: {'Z': -464}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111010; Y = 7'b1111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1083,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b1100001; // Expected: {'Z': -31}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b1100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1084,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100001; Y = 7'b1000110; // Expected: {'Z': 1798}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100001; Y = 7'b1000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1085,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010001; Y = 7'b0011010; // Expected: {'Z': -1222}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010001; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1086,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000111; Y = 7'b0011110; // Expected: {'Z': 210}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000111; Y = 7'b0011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1087,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b1010101; // Expected: {'Z': 1462}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b1010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1088,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000110; Y = 7'b1111010; // Expected: {'Z': -36}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000110; Y = 7'b1111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1089,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111011; Y = 7'b1010100; // Expected: {'Z': -2596}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111011; Y = 7'b1010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1090,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2596
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111010; Y = 7'b1001010; // Expected: {'Z': -3132}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111010; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1091,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110011; Y = 7'b1101000; // Expected: {'Z': -1224}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110011; Y = 7'b1101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1092,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b1100100; // Expected: {'Z': 476}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b1100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1093,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 476
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b1001010; // Expected: {'Z': 2268}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1094,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2268
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b0111100; // Expected: {'Z': -1680}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b0111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1095,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010000; Y = 7'b1010011; // Expected: {'Z': -720}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010000; Y = 7'b1010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1096,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111001; Y = 7'b1001100; // Expected: {'Z': 364}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111001; Y = 7'b1001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1097,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b0110111; // Expected: {'Z': 55}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b0110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1098,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b0001100; // Expected: {'Z': -756}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b0001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1099,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b0101110; // Expected: {'Z': 138}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b0101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1100,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000100; Y = 7'b0000011; // Expected: {'Z': -180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000100; Y = 7'b0000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1101,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b1111110; // Expected: {'Z': -34}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b1111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1102,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011010; Y = 7'b1010001; // Expected: {'Z': 1786}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011010; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1103,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1786
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111111; Y = 7'b0101011; // Expected: {'Z': 2709}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111111; Y = 7'b0101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1104,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2709
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010011; Y = 7'b1011111; // Expected: {'Z': 1485}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010011; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1105,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1485
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000011; Y = 7'b1100101; // Expected: {'Z': 1647}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000011; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1106,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1647
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b1101110; // Expected: {'Z': -162}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b1101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1107,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110011; Y = 7'b0110000; // Expected: {'Z': -624}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110011; Y = 7'b0110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1108,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011111; Y = 7'b0010111; // Expected: {'Z': -759}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011111; Y = 7'b0010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1109,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -759
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b1011100; // Expected: {'Z': -1872}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b1011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1110,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1872
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011010; Y = 7'b0111010; // Expected: {'Z': 1508}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011010; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1111,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1508
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111111; Y = 7'b1111100; // Expected: {'Z': -252}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111111; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1112,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010101; Y = 7'b1000100; // Expected: {'Z': 2580}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010101; Y = 7'b1000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1113,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b1010001; // Expected: {'Z': 1598}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1114,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1598
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b0101011; // Expected: {'Z': -1290}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b0101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1115,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1290
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111100; Y = 7'b1111011; // Expected: {'Z': -300}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111100; Y = 7'b1111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1116,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001000; Y = 7'b1101011; // Expected: {'Z': -168}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001000; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1117,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000111; Y = 7'b1001010; // Expected: {'Z': 3078}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000111; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1118,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3078
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011011; Y = 7'b0011000; // Expected: {'Z': 648}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011011; Y = 7'b0011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1119,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000111; Y = 7'b0010101; // Expected: {'Z': 147}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000111; Y = 7'b0010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1120,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b1110100; // Expected: {'Z': -240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1121,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b1101010; // Expected: {'Z': 66}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b1101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1122,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010000; Y = 7'b1010100; // Expected: {'Z': -704}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010000; Y = 7'b1010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1123,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -704
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b0111111; // Expected: {'Z': -1197}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b0111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1124,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111000; Y = 7'b0101101; // Expected: {'Z': -360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111000; Y = 7'b0101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1125,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110111; Y = 7'b1101011; // Expected: {'Z': 189}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110111; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1126,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010011; Y = 7'b0001110; // Expected: {'Z': 266}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010011; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1127,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 266
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011001; Y = 7'b1000010; // Expected: {'Z': -1550}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011001; Y = 7'b1000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1128,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001100; Y = 7'b1010111; // Expected: {'Z': -492}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001100; Y = 7'b1010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1129,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -492
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010101; Y = 7'b1001101; // Expected: {'Z': 2193}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010101; Y = 7'b1001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1130,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2193
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011001; Y = 7'b0011000; // Expected: {'Z': 600}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011001; Y = 7'b0011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1131,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110011; Y = 7'b1100101; // Expected: {'Z': -1377}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110011; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1132,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1377
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b0101011; // Expected: {'Z': -516}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b0101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1133,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -516
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b0000011; // Expected: {'Z': 186}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b0000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1134,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010111; Y = 7'b0010001; // Expected: {'Z': -697}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010111; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1135,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -697
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000010; Y = 7'b1010011; // Expected: {'Z': -90}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000010; Y = 7'b1010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1136,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111010; Y = 7'b1111001; // Expected: {'Z': -406}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111010; Y = 7'b1111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1137,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -406
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000100; Y = 7'b1000011; // Expected: {'Z': 3660}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000100; Y = 7'b1000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1138,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b1001110; // Expected: {'Z': -450}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b1001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1139,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111011; Y = 7'b1001011; // Expected: {'Z': 265}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111011; Y = 7'b1001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1140,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 265
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b1111101; // Expected: {'Z': 57}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1141,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111101; Y = 7'b0001101; // Expected: {'Z': 793}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111101; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1142,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 793
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100100; Y = 7'b1001111; // Expected: {'Z': -1764}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100100; Y = 7'b1001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1143,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1764
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011011; Y = 7'b1101001; // Expected: {'Z': -621}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011011; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1144,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -621
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b1110001; // Expected: {'Z': 600}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b1110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1145,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011111; Y = 7'b0101010; // Expected: {'Z': -1386}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011111; Y = 7'b0101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1146,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1386
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b0010011; // Expected: {'Z': 380}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b0010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1147,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 380
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111000; Y = 7'b1101001; // Expected: {'Z': 184}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111000; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1148,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b1100101; // Expected: {'Z': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1149,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100100; Y = 7'b1011100; // Expected: {'Z': -1296}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100100; Y = 7'b1011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1150,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110000; Y = 7'b1101111; // Expected: {'Z': -816}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110000; Y = 7'b1101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1151,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110000; Y = 7'b0000110; // Expected: {'Z': 288}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110000; Y = 7'b0000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1152,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101011; Y = 7'b0100010; // Expected: {'Z': -714}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101011; Y = 7'b0100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1153,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -714
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100011; Y = 7'b0011110; // Expected: {'Z': -870}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100011; Y = 7'b0011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1154,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -870
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010011; Y = 7'b0010011; // Expected: {'Z': 361}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010011; Y = 7'b0010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1155,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 361
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110111; Y = 7'b1000100; // Expected: {'Z': -3300}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110111; Y = 7'b1000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1156,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011100; Y = 7'b1100011; // Expected: {'Z': -812}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011100; Y = 7'b1100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1157,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -812
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b1000111; // Expected: {'Z': 684}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b1000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1158,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 684
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011110; Y = 7'b0001110; // Expected: {'Z': 420}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011110; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1159,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110011; Y = 7'b1001101; // Expected: {'Z': -2601}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110011; Y = 7'b1001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1160,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2601
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011011; Y = 7'b0011101; // Expected: {'Z': -1073}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011011; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1161,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1073
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b0010100; // Expected: {'Z': -20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b0010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1162,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b1110010; // Expected: {'Z': -868}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b1110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1163,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -868
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100001; Y = 7'b1011011; // Expected: {'Z': 1147}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100001; Y = 7'b1011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1164,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001101; Y = 7'b1000010; // Expected: {'Z': -806}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001101; Y = 7'b1000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1165,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -806
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000101; Y = 7'b0011111; // Expected: {'Z': 155}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000101; Y = 7'b0011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1166,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b1101110; // Expected: {'Z': 216}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b1101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1167,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000010; Y = 7'b0010110; // Expected: {'Z': -1364}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000010; Y = 7'b0010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1168,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111011; Y = 7'b0100010; // Expected: {'Z': -170}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111011; Y = 7'b0100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1169,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b0111110; // Expected: {'Z': -1116}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b0111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1170,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111100; Y = 7'b1100001; // Expected: {'Z': 124}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111100; Y = 7'b1100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1171,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110010; Y = 7'b0001011; // Expected: {'Z': -154}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110010; Y = 7'b0001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1172,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010111; Y = 7'b0110110; // Expected: {'Z': -2214}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010111; Y = 7'b0110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1173,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001011; Y = 7'b1100101; // Expected: {'Z': -297}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001011; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1174,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -297
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b1000000; // Expected: {'Z': 1280}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b1000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1175,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011001; Y = 7'b0001111; // Expected: {'Z': -585}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011001; Y = 7'b0001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1176,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -585
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b1001010; // Expected: {'Z': -2430}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1177,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b1110100; // Expected: {'Z': 144}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1178,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010111; Y = 7'b0101000; // Expected: {'Z': 920}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010111; Y = 7'b0101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1179,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b1010001; // Expected: {'Z': -423}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1180,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -423
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010100; Y = 7'b1110000; // Expected: {'Z': 704}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010100; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1181,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 704
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011001; Y = 7'b0111011; // Expected: {'Z': -2301}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011001; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1182,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2301
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b1100101; // Expected: {'Z': 756}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1183,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011111; Y = 7'b0110101; // Expected: {'Z': -1749}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011111; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1184,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1749
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010010; Y = 7'b1011110; // Expected: {'Z': -612}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010010; Y = 7'b1011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1185,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b0000011; // Expected: {'Z': 63}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b0000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1186,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000000; Y = 7'b0011101; // Expected: {'Z': -1856}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000000; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1187,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111001; Y = 7'b0111010; // Expected: {'Z': 3306}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111001; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1188,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3306
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b0011000; // Expected: {'Z': -552}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b0011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1189,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b1110101; // Expected: {'Z': -187}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b1110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1190,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011001; Y = 7'b0011100; // Expected: {'Z': -1092}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011001; Y = 7'b0011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1191,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1092
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001101; Y = 7'b0101101; // Expected: {'Z': -2295}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001101; Y = 7'b0101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1192,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2295
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000110; Y = 7'b1110000; // Expected: {'Z': 928}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000110; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1193,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 928
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000010; Y = 7'b1101111; // Expected: {'Z': 1054}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000010; Y = 7'b1101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1194,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1054
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010010; Y = 7'b0100010; // Expected: {'Z': -1564}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010010; Y = 7'b0100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1195,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1564
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101000; Y = 7'b1101101; // Expected: {'Z': 456}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101000; Y = 7'b1101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1196,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100010; Y = 7'b1100010; // Expected: {'Z': -1020}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100010; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1197,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1020
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010000; Y = 7'b0111001; // Expected: {'Z': 912}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010000; Y = 7'b0111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1198,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 912
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b0000010; // Expected: {'Z': -36}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1199,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b1010110; // Expected: {'Z': -2184}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1200,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b0001111; // Expected: {'Z': 360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b0001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1201,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111010; Y = 7'b0000001; // Expected: {'Z': -6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111010; Y = 7'b0000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1202,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001101; Y = 7'b0000111; // Expected: {'Z': 91}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001101; Y = 7'b0000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1203,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011011; Y = 7'b1001001; // Expected: {'Z': 2035}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011011; Y = 7'b1001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1204,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2035
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011100; Y = 7'b0011000; // Expected: {'Z': 672}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011100; Y = 7'b0011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1205,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100111; Y = 7'b1001010; // Expected: {'Z': 1350}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100111; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1206,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111100; Y = 7'b0100101; // Expected: {'Z': 2220}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111100; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1207,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010011; Y = 7'b1000011; // Expected: {'Z': 2745}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010011; Y = 7'b1000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1208,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2745
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001110; Y = 7'b0110100; // Expected: {'Z': 728}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001110; Y = 7'b0110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1209,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010011; Y = 7'b1101100; // Expected: {'Z': -380}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010011; Y = 7'b1101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1210,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -380
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b1000001; // Expected: {'Z': 63}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b1000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1211,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b0010111; // Expected: {'Z': -460}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b0010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1212,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -460
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001101; Y = 7'b0001011; // Expected: {'Z': -561}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001101; Y = 7'b0001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1213,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -561
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111001; Y = 7'b1001100; // Expected: {'Z': -2964}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111001; Y = 7'b1001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1214,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2964
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b0100000; // Expected: {'Z': -1088}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b0100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1215,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1088
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000011; Y = 7'b1010000; // Expected: {'Z': 2928}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000011; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1216,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2928
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101111; Y = 7'b1000110; // Expected: {'Z': -2726}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101111; Y = 7'b1000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1217,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2726
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100011; Y = 7'b1001010; // Expected: {'Z': 1566}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100011; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1218,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1566
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110111; Y = 7'b0111011; // Expected: {'Z': 3245}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110111; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1219,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011010; Y = 7'b1000101; // Expected: {'Z': 2242}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011010; Y = 7'b1000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1220,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111110; Y = 7'b1101000; // Expected: {'Z': 48}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111110; Y = 7'b1101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1221,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101110; Y = 7'b0111000; // Expected: {'Z': 2576}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101110; Y = 7'b0111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1222,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000010; Y = 7'b0010010; // Expected: {'Z': -1116}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000010; Y = 7'b0010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1223,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b0010100; // Expected: {'Z': -640}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b0010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1224,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111001; Y = 7'b0110000; // Expected: {'Z': 2736}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111001; Y = 7'b0110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1225,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000000; Y = 7'b0011011; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000000; Y = 7'b0011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1226,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b0011101; // Expected: {'Z': -1160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1227,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011011; Y = 7'b0001010; // Expected: {'Z': -370}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011011; Y = 7'b0001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1228,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -370
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100001; Y = 7'b0010111; // Expected: {'Z': -713}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100001; Y = 7'b0010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1229,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -713
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101110; Y = 7'b0111000; // Expected: {'Z': 2576}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101110; Y = 7'b0111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1230,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011100; Y = 7'b1000111; // Expected: {'Z': -1596}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011100; Y = 7'b1000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1231,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1596
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b1001110; // Expected: {'Z': -3100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b1001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1232,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100010; Y = 7'b0011101; // Expected: {'Z': 986}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100010; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1233,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 986
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001101; Y = 7'b0011110; // Expected: {'Z': -1530}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001101; Y = 7'b0011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1234,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1530
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101001; Y = 7'b1001011; // Expected: {'Z': -2173}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101001; Y = 7'b1001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1235,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2173
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000011; Y = 7'b0011010; // Expected: {'Z': -1586}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000011; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1236,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1586
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b0001101; // Expected: {'Z': 117}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1237,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b1111011; // Expected: {'Z': -5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b1111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1238,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b0110001; // Expected: {'Z': -490}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b0110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1239,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -490
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001111; Y = 7'b1111010; // Expected: {'Z': 294}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001111; Y = 7'b1111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1240,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 294
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111001; Y = 7'b0111100; // Expected: {'Z': 3420}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111001; Y = 7'b0111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1241,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011101; Y = 7'b1101101; // Expected: {'Z': -551}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011101; Y = 7'b1101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1242,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -551
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000111; Y = 7'b0000110; // Expected: {'Z': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000111; Y = 7'b0000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1243,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000100; Y = 7'b1110000; // Expected: {'Z': -64}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000100; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1244,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110011; Y = 7'b1011111; // Expected: {'Z': 429}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110011; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1245,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 429
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101111; Y = 7'b0101010; // Expected: {'Z': 1974}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101111; Y = 7'b0101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1246,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1974
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b0101111; // Expected: {'Z': -1410}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b0101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1247,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1410
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001111; Y = 7'b1000000; // Expected: {'Z': -960}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001111; Y = 7'b1000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1248,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001111; Y = 7'b1011111; // Expected: {'Z': -495}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001111; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1249,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -495
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b1000111; // Expected: {'Z': 2052}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b1000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1250,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2052
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001010; Y = 7'b0010111; // Expected: {'Z': -1242}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001010; Y = 7'b0010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1251,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101010; Y = 7'b1000101; // Expected: {'Z': -2478}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101010; Y = 7'b1000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1252,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2478
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b0101101; // Expected: {'Z': -1440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b0101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1253,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100010; Y = 7'b1010110; // Expected: {'Z': -1428}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100010; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1254,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1428
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000010; Y = 7'b1100010; // Expected: {'Z': -60}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000010; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1255,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b1110100; // Expected: {'Z': 480}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1256,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100000; Y = 7'b1101110; // Expected: {'Z': -576}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100000; Y = 7'b1101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1257,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001010; Y = 7'b1001000; // Expected: {'Z': -560}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001010; Y = 7'b1001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1258,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b1100000; // Expected: {'Z': 1088}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b1100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1259,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1088
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010001; Y = 7'b0000101; // Expected: {'Z': -235}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010001; Y = 7'b0000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1260,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -235
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b0101000; // Expected: {'Z': 360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b0101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1261,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101011; Y = 7'b0101101; // Expected: {'Z': 1935}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101011; Y = 7'b0101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1262,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1935
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010111; Y = 7'b0101010; // Expected: {'Z': -1722}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010111; Y = 7'b0101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1263,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1722
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111001; Y = 7'b1011001; // Expected: {'Z': 273}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111001; Y = 7'b1011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1264,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 273
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b1110000; // Expected: {'Z': 480}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1265,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b1010110; // Expected: {'Z': 1260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1266,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111011; Y = 7'b0010010; // Expected: {'Z': 1062}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111011; Y = 7'b0010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1267,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1062
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110010; Y = 7'b1000010; // Expected: {'Z': 868}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110010; Y = 7'b1000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1268,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 868
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b0110101; // Expected: {'Z': 2385}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1269,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2385
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b1101000; // Expected: {'Z': -576}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b1101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1270,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001011; Y = 7'b0000001; // Expected: {'Z': -53}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001011; Y = 7'b0000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1271,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b0011101; // Expected: {'Z': 1537}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1272,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1537
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b0101101; // Expected: {'Z': 900}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b0101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1273,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001100; Y = 7'b0101111; // Expected: {'Z': 564}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001100; Y = 7'b0101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1274,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 564
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011111; Y = 7'b0010000; // Expected: {'Z': 496}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011111; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1275,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011010; Y = 7'b0001000; // Expected: {'Z': -304}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011010; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1276,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -304
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100101; Y = 7'b0100001; // Expected: {'Z': 1221}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100101; Y = 7'b0100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1277,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000000; Y = 7'b0011010; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000000; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1278,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010110; Y = 7'b0010110; // Expected: {'Z': 484}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010110; Y = 7'b0010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1279,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 484
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000100; Y = 7'b0111001; // Expected: {'Z': 228}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000100; Y = 7'b0111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1280,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101110; Y = 7'b1010001; // Expected: {'Z': -2162}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101110; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1281,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001100; Y = 7'b0010011; // Expected: {'Z': -988}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001100; Y = 7'b0010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1282,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -988
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b0001100; // Expected: {'Z': 288}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b0001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1283,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011100; Y = 7'b1001000; // Expected: {'Z': -1568}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011100; Y = 7'b1001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1284,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1568
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010011; Y = 7'b1110100; // Expected: {'Z': 540}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010011; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1285,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000011; Y = 7'b1001111; // Expected: {'Z': 2989}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000011; Y = 7'b1001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1286,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2989
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100100; Y = 7'b0000100; // Expected: {'Z': 144}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100100; Y = 7'b0000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1287,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000111; Y = 7'b1000011; // Expected: {'Z': 3477}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000111; Y = 7'b1000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1288,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3477
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000110; Y = 7'b1000111; // Expected: {'Z': 3306}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000110; Y = 7'b1000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1289,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3306
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101010; Y = 7'b0100100; // Expected: {'Z': -792}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101010; Y = 7'b0100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1290,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b1101101; // Expected: {'Z': -1007}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b1101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1291,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1007
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010111; Y = 7'b0110001; // Expected: {'Z': -2009}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010111; Y = 7'b0110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1292,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2009
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100001; Y = 7'b1101011; // Expected: {'Z': -693}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100001; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1293,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -693
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b0101000; // Expected: {'Z': 2480}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b0101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1294,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000010; Y = 7'b1010000; // Expected: {'Z': -96}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000010; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1295,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010011; Y = 7'b0110010; // Expected: {'Z': -2250}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010011; Y = 7'b0110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1296,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b0101001; // Expected: {'Z': -410}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1297,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -410
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b1011011; // Expected: {'Z': 1480}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b1011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1298,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b1001011; // Expected: {'Z': 1219}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b1001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1299,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1219
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011010; Y = 7'b0111011; // Expected: {'Z': 1534}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011010; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1300,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1534
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101010; Y = 7'b1100000; // Expected: {'Z': -1344}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101010; Y = 7'b1100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1301,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1344
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101100; Y = 7'b0110011; // Expected: {'Z': 2244}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101100; Y = 7'b0110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1302,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101110; Y = 7'b1110100; // Expected: {'Z': -552}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101110; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1303,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b0011001; // Expected: {'Z': 425}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b0011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1304,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 425
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001100; Y = 7'b0001101; // Expected: {'Z': 156}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001100; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1305,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001110; Y = 7'b0110110; // Expected: {'Z': 756}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001110; Y = 7'b0110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1306,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101011; Y = 7'b1111100; // Expected: {'Z': 84}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101011; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1307,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b1100110; // Expected: {'Z': 728}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b1100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1308,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b0000100; // Expected: {'Z': -120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b0000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1309,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b1001110; // Expected: {'Z': -3100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b1001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1310,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100110; Y = 7'b0111111; // Expected: {'Z': 2394}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100110; Y = 7'b0111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1311,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2394
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011011; Y = 7'b0011101; // Expected: {'Z': -1073}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011011; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1312,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1073
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101000; Y = 7'b0000100; // Expected: {'Z': -96}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101000; Y = 7'b0000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1313,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001010; Y = 7'b0100000; // Expected: {'Z': -1728}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001010; Y = 7'b0100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1314,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b0011110; // Expected: {'Z': -1440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b0011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1315,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b0101101; // Expected: {'Z': -855}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b0101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1316,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -855
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000011; Y = 7'b0111011; // Expected: {'Z': -3599}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000011; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1317,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3599
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b1010100; // Expected: {'Z': 2772}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b1010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1318,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2772
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111001; Y = 7'b1111110; // Expected: {'Z': -114}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111001; Y = 7'b1111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1319,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101011; Y = 7'b1100100; // Expected: {'Z': -1204}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101011; Y = 7'b1100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1320,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100101; Y = 7'b1100000; // Expected: {'Z': 864}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100101; Y = 7'b1100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1321,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 864
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b0010110; // Expected: {'Z': -66}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b0010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1322,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010011; Y = 7'b1101000; // Expected: {'Z': -456}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010011; Y = 7'b1101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1323,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001101; Y = 7'b0100011; // Expected: {'Z': -1785}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001101; Y = 7'b0100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1324,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1785
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100001; Y = 7'b0001001; // Expected: {'Z': -279}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100001; Y = 7'b0001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1325,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -279
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000101; Y = 7'b1001100; // Expected: {'Z': 3068}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000101; Y = 7'b1001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1326,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3068
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101001; Y = 7'b1000011; // Expected: {'Z': -2501}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101001; Y = 7'b1000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1327,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2501
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100110; Y = 7'b0111011; // Expected: {'Z': 2242}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100110; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1328,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b1110110; // Expected: {'Z': -170}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1329,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b0101010; // Expected: {'Z': -1344}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b0101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1330,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1344
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b1010111; // Expected: {'Z': -2132}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b1010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1331,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100001; Y = 7'b1101100; // Expected: {'Z': 620}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100001; Y = 7'b1101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1332,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010000; Y = 7'b1001101; // Expected: {'Z': -816}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010000; Y = 7'b1001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1333,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011101; Y = 7'b1011100; // Expected: {'Z': 1260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011101; Y = 7'b1011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1334,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b1100110; // Expected: {'Z': 1248}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b1100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1335,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010011; Y = 7'b0101001; // Expected: {'Z': 779}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010011; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1336,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 779
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b1010110; // Expected: {'Z': 966}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1337,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 966
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110000; Y = 7'b0101111; // Expected: {'Z': 2256}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110000; Y = 7'b0101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1338,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2256
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101111; Y = 7'b1100110; // Expected: {'Z': -1222}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101111; Y = 7'b1100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1339,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010100; Y = 7'b0101100; // Expected: {'Z': -1936}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010100; Y = 7'b0101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1340,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1936
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b0011110; // Expected: {'Z': -1260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b0011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1341,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010001; Y = 7'b1011000; // Expected: {'Z': 1880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010001; Y = 7'b1011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1342,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100101; Y = 7'b0101010; // Expected: {'Z': -1134}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100101; Y = 7'b0101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1343,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001001; Y = 7'b0010100; // Expected: {'Z': -1100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001001; Y = 7'b0010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1344,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111000; Y = 7'b0011011; // Expected: {'Z': 1512}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111000; Y = 7'b0011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1345,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1512
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110111; Y = 7'b1100010; // Expected: {'Z': 270}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110111; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1346,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 270
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011001; Y = 7'b1011011; // Expected: {'Z': 1443}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011001; Y = 7'b1011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1347,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1443
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101011; Y = 7'b1010101; // Expected: {'Z': -1849}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101011; Y = 7'b1010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1348,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1849
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b1101000; // Expected: {'Z': 816}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b1101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1349,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111111; Y = 7'b1110110; // Expected: {'Z': -630}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111111; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1350,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -630
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001101; Y = 7'b0111100; // Expected: {'Z': 780}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001101; Y = 7'b0111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1351,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b0101001; // Expected: {'Z': 1845}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1352,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1845
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111111; Y = 7'b1000101; // Expected: {'Z': -3717}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111111; Y = 7'b1000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1353,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3717
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b0111011; // Expected: {'Z': -1652}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1354,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1652
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000010; Y = 7'b1011000; // Expected: {'Z': -80}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000010; Y = 7'b1011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1355,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001010; Y = 7'b0011011; // Expected: {'Z': 270}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001010; Y = 7'b0011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1356,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 270
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100101; Y = 7'b0101001; // Expected: {'Z': -1107}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100101; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1357,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000111; Y = 7'b1011010; // Expected: {'Z': 2166}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000111; Y = 7'b1011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1358,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001101; Y = 7'b1101101; // Expected: {'Z': 969}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001101; Y = 7'b1101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1359,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 969
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b0010111; // Expected: {'Z': -23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b0010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1360,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b0000101; // Expected: {'Z': -180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b0000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1361,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b0101000; // Expected: {'Z': 2480}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b0101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1362,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b1110011; // Expected: {'Z': -13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1363,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010011; Y = 7'b1001101; // Expected: {'Z': 2295}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010011; Y = 7'b1001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1364,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2295
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110010; Y = 7'b1011111; // Expected: {'Z': -1650}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110010; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1365,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101100; Y = 7'b1001100; // Expected: {'Z': -2288}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101100; Y = 7'b1001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1366,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010000; Y = 7'b0100100; // Expected: {'Z': 576}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010000; Y = 7'b0100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1367,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100110; Y = 7'b1101011; // Expected: {'Z': 546}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100110; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1368,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b0111110; // Expected: {'Z': -1240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b0111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1369,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000100; Y = 7'b1100011; // Expected: {'Z': -116}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000100; Y = 7'b1100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1370,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001100; Y = 7'b1111100; // Expected: {'Z': 208}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001100; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1371,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b1001000; // Expected: {'Z': 672}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b1001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1372,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000000; Y = 7'b0000101; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000000; Y = 7'b0000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1373,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b1011001; // Expected: {'Z': 780}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b1011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1374,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101001; Y = 7'b1110101; // Expected: {'Z': -451}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101001; Y = 7'b1110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1375,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -451
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010111; Y = 7'b1001000; // Expected: {'Z': -1288}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010111; Y = 7'b1001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1376,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000011; Y = 7'b0101001; // Expected: {'Z': -2501}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000011; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1377,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2501
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011011; Y = 7'b1011011; // Expected: {'Z': 1369}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011011; Y = 7'b1011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1378,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1369
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110110; Y = 7'b1110101; // Expected: {'Z': -594}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110110; Y = 7'b1110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1379,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -594
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110010; Y = 7'b1010111; // Expected: {'Z': 574}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110010; Y = 7'b1010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1380,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 574
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111111; Y = 7'b0110010; // Expected: {'Z': 3150}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111111; Y = 7'b0110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1381,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010101; Y = 7'b0011010; // Expected: {'Z': -1118}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010101; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1382,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010111; Y = 7'b1000000; // Expected: {'Z': -1472}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010111; Y = 7'b1000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1383,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1472
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111010; Y = 7'b0100111; // Expected: {'Z': -234}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111010; Y = 7'b0100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1384,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010010; Y = 7'b0001010; // Expected: {'Z': -460}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010010; Y = 7'b0001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1385,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -460
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101001; Y = 7'b0111000; // Expected: {'Z': 2296}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101001; Y = 7'b0111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1386,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000101; Y = 7'b0101001; // Expected: {'Z': -2419}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000101; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1387,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2419
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110111; Y = 7'b1101001; // Expected: {'Z': 207}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110111; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1388,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 207
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b1110011; // Expected: {'Z': 156}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1389,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111110; Y = 7'b1101010; // Expected: {'Z': 44}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111110; Y = 7'b1101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1390,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100100; Y = 7'b1010010; // Expected: {'Z': -1656}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100100; Y = 7'b1010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1391,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1656
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111100; Y = 7'b0010001; // Expected: {'Z': -68}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111100; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1392,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000110; Y = 7'b0000011; // Expected: {'Z': -174}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000110; Y = 7'b0000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1393,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010011; Y = 7'b1001100; // Expected: {'Z': -988}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010011; Y = 7'b1001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1394,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -988
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111110; Y = 7'b0001010; // Expected: {'Z': -20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111110; Y = 7'b0001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1395,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000110; Y = 7'b1010000; // Expected: {'Z': -288}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000110; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1396,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100110; Y = 7'b1101111; // Expected: {'Z': 442}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100110; Y = 7'b1101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1397,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 442
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111011; Y = 7'b0000110; // Expected: {'Z': 354}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111011; Y = 7'b0000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1398,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 354
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010100; Y = 7'b1101100; // Expected: {'Z': 880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010100; Y = 7'b1101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1399,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b0111000; // Expected: {'Z': -2352}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b0111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1400,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001101; Y = 7'b0111100; // Expected: {'Z': -3060}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001101; Y = 7'b0111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1401,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001111; Y = 7'b1100101; // Expected: {'Z': 1323}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001111; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1402,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1323
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101011; Y = 7'b1011011; // Expected: {'Z': 777}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101011; Y = 7'b1011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1403,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 777
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b1100110; // Expected: {'Z': 1092}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b1100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1404,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1092
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100101; Y = 7'b0111110; // Expected: {'Z': -1674}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100101; Y = 7'b0111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1405,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1674
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100111; Y = 7'b1000111; // Expected: {'Z': 1425}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100111; Y = 7'b1000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1406,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1425
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001101; Y = 7'b0101110; // Expected: {'Z': 598}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001101; Y = 7'b0101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1407,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 598
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001111; Y = 7'b0001111; // Expected: {'Z': 225}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001111; Y = 7'b0001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1408,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000000; Y = 7'b0010110; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000000; Y = 7'b0010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1409,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010110; Y = 7'b0110111; // Expected: {'Z': 1210}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010110; Y = 7'b0110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1410,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101011; Y = 7'b0100111; // Expected: {'Z': 1677}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101011; Y = 7'b0100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1411,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1677
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b1100010; // Expected: {'Z': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1412,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111011; Y = 7'b1010110; // Expected: {'Z': -2478}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111011; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1413,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2478
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b1101111; // Expected: {'Z': 51}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b1101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1414,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b0010100; // Expected: {'Z': -200}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b0010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1415,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100111; Y = 7'b0100010; // Expected: {'Z': 1326}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100111; Y = 7'b0100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1416,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1326
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111110; Y = 7'b1100101; // Expected: {'Z': 54}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111110; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1417,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b0100111; // Expected: {'Z': 2028}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b0100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1418,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2028
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100101; Y = 7'b1011000; // Expected: {'Z': -1480}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100101; Y = 7'b1011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1419,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b0000111; // Expected: {'Z': -294}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b0000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1420,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -294
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100110; Y = 7'b1110000; // Expected: {'Z': 416}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100110; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1421,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001010; Y = 7'b1101100; // Expected: {'Z': -200}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001010; Y = 7'b1101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1422,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011010; Y = 7'b0011110; // Expected: {'Z': 780}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011010; Y = 7'b0011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1423,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b1110100; // Expected: {'Z': -252}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1424,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111011; Y = 7'b0011000; // Expected: {'Z': -120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111011; Y = 7'b0011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1425,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b0001111; // Expected: {'Z': -150}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b0001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1426,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010000; Y = 7'b0111010; // Expected: {'Z': 928}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010000; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1427,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 928
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010101; Y = 7'b0111011; // Expected: {'Z': -2537}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010101; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1428,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2537
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b0010011; // Expected: {'Z': -342}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b0010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1429,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -342
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010111; Y = 7'b0000110; // Expected: {'Z': -246}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010111; Y = 7'b0000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1430,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b1010111; // Expected: {'Z': 1968}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b1010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1431,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1968
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110110; Y = 7'b1000110; // Expected: {'Z': -3132}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110110; Y = 7'b1000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1432,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110111; Y = 7'b0111011; // Expected: {'Z': -531}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110111; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1433,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -531
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b1100101; // Expected: {'Z': 810}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1434,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 810
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000110; Y = 7'b0101110; // Expected: {'Z': -2668}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000110; Y = 7'b0101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1435,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2668
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000100; Y = 7'b1111110; // Expected: {'Z': 120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000100; Y = 7'b1111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1436,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b0100011; // Expected: {'Z': 1855}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b0100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1437,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1855
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000110; Y = 7'b1100101; // Expected: {'Z': -162}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000110; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1438,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101010; Y = 7'b0000100; // Expected: {'Z': -88}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101010; Y = 7'b0000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1439,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101000; Y = 7'b1111001; // Expected: {'Z': -280}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101000; Y = 7'b1111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1440,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000000; Y = 7'b1010001; // Expected: {'Z': 3008}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000000; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1441,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111000; Y = 7'b0101111; // Expected: {'Z': -376}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111000; Y = 7'b0101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1442,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -376
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b1011101; // Expected: {'Z': 525}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b1011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1443,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 525
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010011; Y = 7'b1011000; // Expected: {'Z': -760}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010011; Y = 7'b1011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1444,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100001; Y = 7'b1111001; // Expected: {'Z': 217}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100001; Y = 7'b1111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1445,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001101; Y = 7'b1100111; // Expected: {'Z': 1275}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001101; Y = 7'b1100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1446,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1275
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011001; Y = 7'b1001001; // Expected: {'Z': 2145}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011001; Y = 7'b1001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1447,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001110; Y = 7'b1111011; // Expected: {'Z': 250}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001110; Y = 7'b1111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1448,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100100; Y = 7'b1110110; // Expected: {'Z': -360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100100; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1449,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001011; Y = 7'b0111011; // Expected: {'Z': 649}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001011; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1450,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 649
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001111; Y = 7'b0011101; // Expected: {'Z': -1421}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001111; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1451,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1421
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b0101101; // Expected: {'Z': -1350}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b0101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1452,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011011; Y = 7'b0000110; // Expected: {'Z': 162}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011011; Y = 7'b0000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1453,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000110; Y = 7'b0111110; // Expected: {'Z': 372}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000110; Y = 7'b0111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1454,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 372
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010100; Y = 7'b1101011; // Expected: {'Z': 924}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010100; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1455,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 924
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101110; Y = 7'b1001100; // Expected: {'Z': -2392}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101110; Y = 7'b1001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1456,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010011; Y = 7'b0001000; // Expected: {'Z': 152}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010011; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1457,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b0111110; // Expected: {'Z': -186}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b0111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1458,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010101; Y = 7'b0110000; // Expected: {'Z': -2064}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010101; Y = 7'b0110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1459,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2064
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000110; Y = 7'b0100110; // Expected: {'Z': 228}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000110; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1460,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100110; Y = 7'b1010000; // Expected: {'Z': -1824}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100110; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1461,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1824
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011010; Y = 7'b0101000; // Expected: {'Z': -1520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011010; Y = 7'b0101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1462,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b1000001; // Expected: {'Z': 3969}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b1000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1463,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3969
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111100; Y = 7'b1111001; // Expected: {'Z': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111100; Y = 7'b1111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1464,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b0000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b0000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1465,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b1001011; // Expected: {'Z': 2226}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b1001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1466,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2226
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101001; Y = 7'b0010001; // Expected: {'Z': 697}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101001; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1467,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 697
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111011; Y = 7'b0111100; // Expected: {'Z': -300}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111011; Y = 7'b0111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1468,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110110; Y = 7'b1000001; // Expected: {'Z': -3402}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110110; Y = 7'b1000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1469,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3402
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001010; Y = 7'b1110011; // Expected: {'Z': -130}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001010; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1470,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000101; Y = 7'b1010011; // Expected: {'Z': 2655}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000101; Y = 7'b1010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1471,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2655
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100011; Y = 7'b0101011; // Expected: {'Z': 1505}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100011; Y = 7'b0101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1472,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1505
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b0000011; // Expected: {'Z': -51}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b0000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1473,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b0000110; // Expected: {'Z': -60}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b0000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1474,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b1101111; // Expected: {'Z': 544}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b1101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1475,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 544
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001101; Y = 7'b1010101; // Expected: {'Z': -559}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001101; Y = 7'b1010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1476,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -559
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000101; Y = 7'b1110010; // Expected: {'Z': 826}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000101; Y = 7'b1110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1477,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 826
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b1110110; // Expected: {'Z': 120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1478,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b1111110; // Expected: {'Z': -124}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b1111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1479,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b0011100; // Expected: {'Z': -420}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b0011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1480,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b0011011; // Expected: {'Z': -864}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b0011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1481,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -864
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011111; Y = 7'b0101011; // Expected: {'Z': -1419}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011111; Y = 7'b0101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1482,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1419
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000100; Y = 7'b1010001; // Expected: {'Z': -188}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000100; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1483,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111100; Y = 7'b0011110; // Expected: {'Z': 1800}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111100; Y = 7'b0011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1484,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b0011010; // Expected: {'Z': 520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1485,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111101; Y = 7'b0100100; // Expected: {'Z': 2196}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111101; Y = 7'b0100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1486,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010010; Y = 7'b0010010; // Expected: {'Z': -828}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010010; Y = 7'b0010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1487,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010010; Y = 7'b0001100; // Expected: {'Z': -552}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010010; Y = 7'b0001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1488,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001111; Y = 7'b1001010; // Expected: {'Z': 2646}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001111; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1489,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2646
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101010; Y = 7'b0000010; // Expected: {'Z': -44}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101010; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1490,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100000; Y = 7'b1111111; // Expected: {'Z': -32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100000; Y = 7'b1111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1491,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b0011110; // Expected: {'Z': 1860}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b0011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1492,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1860
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111000; Y = 7'b1110110; // Expected: {'Z': -560}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111000; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1493,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000100; Y = 7'b1110001; // Expected: {'Z': -60}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000100; Y = 7'b1110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1494,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b1110000; // Expected: {'Z': 448}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1495,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 448
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000010; Y = 7'b1110100; // Expected: {'Z': 744}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000010; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1496,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 744
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001100; Y = 7'b1011100; // Expected: {'Z': 1872}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001100; Y = 7'b1011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1497,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1872
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101000; Y = 7'b0111100; // Expected: {'Z': -1440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101000; Y = 7'b0111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1498,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101010; Y = 7'b1110100; // Expected: {'Z': -504}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101010; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1499,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110001; Y = 7'b0101100; // Expected: {'Z': 2156}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110001; Y = 7'b0101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1500,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001111; Y = 7'b1010100; // Expected: {'Z': 2156}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001111; Y = 7'b1010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1501,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b1000110; // Expected: {'Z': 986}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b1000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1502,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 986
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011011; Y = 7'b1000110; // Expected: {'Z': 2146}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011011; Y = 7'b1000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1503,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100001; Y = 7'b1111100; // Expected: {'Z': 124}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100001; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1504,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b0001010; // Expected: {'Z': -10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b0001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1505,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b1111011; // Expected: {'Z': -85}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b1111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1506,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -85
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001100; Y = 7'b0001100; // Expected: {'Z': -624}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001100; Y = 7'b0001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1507,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011111; Y = 7'b1111100; // Expected: {'Z': -124}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011111; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1508,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b1011010; // Expected: {'Z': -2014}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b1011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1509,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2014
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b1000111; // Expected: {'Z': 969}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b1000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1510,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 969
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b0010110; // Expected: {'Z': 1364}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b0010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1511,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111101; Y = 7'b0111011; // Expected: {'Z': 3599}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111101; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1512,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3599
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b1110011; // Expected: {'Z': -39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1513,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000010; Y = 7'b0110010; // Expected: {'Z': -3100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000010; Y = 7'b0110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1514,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100011; Y = 7'b1000111; // Expected: {'Z': 1653}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100011; Y = 7'b1000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1515,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1653
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110000; Y = 7'b1111100; // Expected: {'Z': 64}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110000; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1516,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011100; Y = 7'b1000010; // Expected: {'Z': -1736}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011100; Y = 7'b1000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1517,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b1100110; // Expected: {'Z': -624}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b1100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1518,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b1100100; // Expected: {'Z': -672}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b1100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1519,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001010; Y = 7'b0111000; // Expected: {'Z': 560}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001010; Y = 7'b0111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1520,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000010; Y = 7'b1001011; // Expected: {'Z': -106}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000010; Y = 7'b1001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1521,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b1010000; // Expected: {'Z': -2544}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1522,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2544
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b0010111; // Expected: {'Z': -345}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b0010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1523,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -345
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101001; Y = 7'b1111101; // Expected: {'Z': -123}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101001; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1524,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -123
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000110; Y = 7'b1101010; // Expected: {'Z': -132}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000110; Y = 7'b1101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1525,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b0011110; // Expected: {'Z': 1590}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b0011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1526,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1590
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b0010010; // Expected: {'Z': -18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b0010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1527,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001010; Y = 7'b0001110; // Expected: {'Z': -756}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001010; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1528,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000110; Y = 7'b1001111; // Expected: {'Z': 2842}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000110; Y = 7'b1001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1529,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2842
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b1100011; // Expected: {'Z': -609}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b1100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1530,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -609
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010010; Y = 7'b0101111; // Expected: {'Z': -2162}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010010; Y = 7'b0101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1531,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b0010101; // Expected: {'Z': 1113}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b0010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1532,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101010; Y = 7'b1100001; // Expected: {'Z': -1302}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101010; Y = 7'b1100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1533,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1302
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010001; Y = 7'b1000010; // Expected: {'Z': 2914}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010001; Y = 7'b1000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1534,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2914
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111111; Y = 7'b1110111; // Expected: {'Z': -567}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111111; Y = 7'b1110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1535,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -567
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b1011100; // Expected: {'Z': 720}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b1011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1536,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011011; Y = 7'b0000111; // Expected: {'Z': -259}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011011; Y = 7'b0000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1537,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -259
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110011; Y = 7'b0000100; // Expected: {'Z': 204}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110011; Y = 7'b0000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1538,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b0001000; // Expected: {'Z': 496}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1539,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001001; Y = 7'b0000001; // Expected: {'Z': -55}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001001; Y = 7'b0000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1540,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110000; Y = 7'b0110001; // Expected: {'Z': -784}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110000; Y = 7'b0110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1541,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101000; Y = 7'b1110011; // Expected: {'Z': 312}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101000; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1542,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 312
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110010; Y = 7'b0110000; // Expected: {'Z': 2400}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110010; Y = 7'b0110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1543,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b1011110; // Expected: {'Z': 1224}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b1011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1544,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111100; Y = 7'b1111110; // Expected: {'Z': -120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111100; Y = 7'b1111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1545,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b1000101; // Expected: {'Z': 1888}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b1000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1546,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110000; Y = 7'b0100101; // Expected: {'Z': 1776}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110000; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1547,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1776
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101110; Y = 7'b1010110; // Expected: {'Z': -1932}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101110; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1548,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1932
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b0000110; // Expected: {'Z': 270}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b0000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1549,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 270
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111011; Y = 7'b0000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111011; Y = 7'b0000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1550,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011111; Y = 7'b1000111; // Expected: {'Z': -1767}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011111; Y = 7'b1000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1551,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1767
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100110; Y = 7'b1111101; // Expected: {'Z': -114}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100110; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1552,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b0001000; // Expected: {'Z': -8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1553,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b0010000; // Expected: {'Z': -320}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1554,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011001; Y = 7'b0000110; // Expected: {'Z': 150}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011001; Y = 7'b0000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1555,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010010; Y = 7'b0001011; // Expected: {'Z': 198}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010010; Y = 7'b0001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1556,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110011; Y = 7'b0100001; // Expected: {'Z': -429}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110011; Y = 7'b0100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1557,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -429
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b0011010; // Expected: {'Z': -26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1558,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101011; Y = 7'b0010110; // Expected: {'Z': 946}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101011; Y = 7'b0010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1559,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 946
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100000; Y = 7'b0100100; // Expected: {'Z': 1152}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100000; Y = 7'b0100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1560,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b1011101; // Expected: {'Z': 1400}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b1011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1561,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100111; Y = 7'b1010011; // Expected: {'Z': 1125}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100111; Y = 7'b1010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1562,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000010; Y = 7'b1010001; // Expected: {'Z': -94}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000010; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1563,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b1011001; // Expected: {'Z': 2457}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b1011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1564,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2457
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000000; Y = 7'b1110011; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000000; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1565,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b1001101; // Expected: {'Z': 765}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b1001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1566,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 765
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b0010001; // Expected: {'Z': -51}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1567,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100010; Y = 7'b0010100; // Expected: {'Z': 680}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100010; Y = 7'b0010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1568,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010000; Y = 7'b0101011; // Expected: {'Z': 688}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010000; Y = 7'b0101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1569,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 688
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001110; Y = 7'b0100110; // Expected: {'Z': -1900}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001110; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1570,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111110; Y = 7'b1011100; // Expected: {'Z': 72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111110; Y = 7'b1011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1571,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000110; Y = 7'b1000000; // Expected: {'Z': -384}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000110; Y = 7'b1000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1572,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -384
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011100; Y = 7'b0101011; // Expected: {'Z': 1204}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011100; Y = 7'b0101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1573,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b1100010; // Expected: {'Z': 690}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1574,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 690
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001110; Y = 7'b0110010; // Expected: {'Z': -2500}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001110; Y = 7'b0110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1575,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001000; Y = 7'b1001101; // Expected: {'Z': 2856}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001000; Y = 7'b1001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1576,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001101; Y = 7'b1111000; // Expected: {'Z': 408}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001101; Y = 7'b1111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1577,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011111; Y = 7'b1000001; // Expected: {'Z': -1953}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011111; Y = 7'b1000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1578,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1953
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110111; Y = 7'b1111001; // Expected: {'Z': 63}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110111; Y = 7'b1111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1579,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b0000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b0000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1580,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010111; Y = 7'b0001100; // Expected: {'Z': -492}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010111; Y = 7'b0001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1581,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -492
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b0010111; // Expected: {'Z': -230}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b0010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1582,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000000; Y = 7'b0111101; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000000; Y = 7'b0111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1583,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b0001011; // Expected: {'Z': 583}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b0001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1584,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 583
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111101; Y = 7'b0010010; // Expected: {'Z': 1098}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111101; Y = 7'b0010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1585,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1098
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b1111000; // Expected: {'Z': -496}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b1111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1586,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100110; Y = 7'b0101110; // Expected: {'Z': 1748}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100110; Y = 7'b0101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1587,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1748
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b0110001; // Expected: {'Z': -3087}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b0110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1588,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3087
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b1001111; // Expected: {'Z': 1127}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b1001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1589,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1127
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b1100101; // Expected: {'Z': 864}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1590,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 864
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b0001100; // Expected: {'Z': -228}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b0001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1591,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110010; Y = 7'b1010110; // Expected: {'Z': -2100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110010; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1592,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010000; Y = 7'b1000110; // Expected: {'Z': -928}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010000; Y = 7'b1000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1593,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -928
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001111; Y = 7'b1001010; // Expected: {'Z': -810}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001111; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1594,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -810
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110101; Y = 7'b0101010; // Expected: {'Z': -462}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110101; Y = 7'b0101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1595,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b1011110; // Expected: {'Z': 408}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b1011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1596,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110111; Y = 7'b1010111; // Expected: {'Z': -2255}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110111; Y = 7'b1010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1597,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b0100001; // Expected: {'Z': 1716}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b0100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1598,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1716
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001010; Y = 7'b0011111; // Expected: {'Z': 310}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001010; Y = 7'b0011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1599,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 310
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011101; Y = 7'b0011100; // Expected: {'Z': -980}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011101; Y = 7'b0011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1600,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101010; Y = 7'b1010100; // Expected: {'Z': 968}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101010; Y = 7'b1010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1601,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 968
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000011; Y = 7'b0110100; // Expected: {'Z': -3172}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000011; Y = 7'b0110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1602,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b1110000; // Expected: {'Z': 544}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1603,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 544
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b0010010; // Expected: {'Z': -648}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b0010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1604,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011011; Y = 7'b0101101; // Expected: {'Z': -1665}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011011; Y = 7'b0101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1605,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1665
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100011; Y = 7'b1111111; // Expected: {'Z': -35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100011; Y = 7'b1111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1606,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b1100111; // Expected: {'Z': 575}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b1100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1607,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 575
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001111; Y = 7'b1100000; // Expected: {'Z': -480}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001111; Y = 7'b1100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1608,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111010; Y = 7'b1100110; // Expected: {'Z': -1508}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111010; Y = 7'b1100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1609,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1508
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111010; Y = 7'b1010100; // Expected: {'Z': 264}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111010; Y = 7'b1010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1610,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010111; Y = 7'b0001010; // Expected: {'Z': -410}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010111; Y = 7'b0001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1611,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -410
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011111; Y = 7'b0011010; // Expected: {'Z': 806}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011111; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1612,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 806
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001100; Y = 7'b0001000; // Expected: {'Z': 96}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001100; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1613,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111000; Y = 7'b1010010; // Expected: {'Z': -2576}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111000; Y = 7'b1010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1614,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b0000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b0000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1615,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100011; Y = 7'b0011010; // Expected: {'Z': 910}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100011; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1616,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 910
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011101; Y = 7'b1111100; // Expected: {'Z': 140}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011101; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1617,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111010; Y = 7'b0111011; // Expected: {'Z': -354}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111010; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1618,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -354
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101011; Y = 7'b0101011; // Expected: {'Z': 1849}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101011; Y = 7'b0101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1619,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1849
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b0101101; // Expected: {'Z': 1080}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b0101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1620,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b0101011; // Expected: {'Z': -731}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b0101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1621,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -731
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b1010100; // Expected: {'Z': 880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b1010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1622,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b0110100; // Expected: {'Z': -1456}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b0110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1623,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100100; Y = 7'b1000001; // Expected: {'Z': -2268}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100100; Y = 7'b1000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1624,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2268
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b0000111; // Expected: {'Z': 147}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b0000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1625,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b0101010; // Expected: {'Z': 882}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b0101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1626,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 882
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100111; Y = 7'b1100010; // Expected: {'Z': -1170}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100111; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1627,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b1101100; // Expected: {'Z': -1040}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b1101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1628,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b1111001; // Expected: {'Z': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b1111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1629,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001101; Y = 7'b1011010; // Expected: {'Z': 1938}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001101; Y = 7'b1011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1630,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1938
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101011; Y = 7'b1010000; // Expected: {'Z': 1008}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101011; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1631,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100100; Y = 7'b0001101; // Expected: {'Z': 468}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100100; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1632,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 468
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b0011000; // Expected: {'Z': -1008}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b0011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1633,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101011; Y = 7'b0111101; // Expected: {'Z': -1281}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101011; Y = 7'b0111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1634,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1281
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b0110000; // Expected: {'Z': -1728}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b0110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1635,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b0101100; // Expected: {'Z': -2112}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b0101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1636,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010100; Y = 7'b1101011; // Expected: {'Z': 924}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010100; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1637,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 924
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011011; Y = 7'b1001010; // Expected: {'Z': -1458}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011011; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1638,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1458
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111111; Y = 7'b0100100; // Expected: {'Z': 2268}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111111; Y = 7'b0100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1639,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2268
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100000; Y = 7'b0111011; // Expected: {'Z': 1888}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100000; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1640,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010110; Y = 7'b1110101; // Expected: {'Z': -242}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010110; Y = 7'b1110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1641,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b1011011; // Expected: {'Z': -111}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b1011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1642,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -111
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100001; Y = 7'b1110111; // Expected: {'Z': 279}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100001; Y = 7'b1110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1643,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 279
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001011; Y = 7'b1101111; // Expected: {'Z': -187}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001011; Y = 7'b1101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1644,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b0100000; // Expected: {'Z': 640}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b0100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1645,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b1010010; // Expected: {'Z': 1564}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b1010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1646,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1564
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001011; Y = 7'b0110000; // Expected: {'Z': 528}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001011; Y = 7'b0110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1647,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111000; Y = 7'b0010100; // Expected: {'Z': -160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111000; Y = 7'b0010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1648,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001010; Y = 7'b1110100; // Expected: {'Z': 648}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001010; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1649,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101010; Y = 7'b0011000; // Expected: {'Z': -528}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101010; Y = 7'b0011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1650,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111110; Y = 7'b1101100; // Expected: {'Z': 40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111110; Y = 7'b1101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1651,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111001; Y = 7'b1110010; // Expected: {'Z': -798}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111001; Y = 7'b1110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1652,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101110; Y = 7'b0010111; // Expected: {'Z': 1058}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101110; Y = 7'b0010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1653,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1058
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b0010111; // Expected: {'Z': -437}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b0010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1654,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -437
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000111; Y = 7'b0000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000111; Y = 7'b0000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1655,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111100; Y = 7'b0011111; // Expected: {'Z': 1860}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111100; Y = 7'b0011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1656,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1860
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111100; Y = 7'b0001110; // Expected: {'Z': 840}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111100; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1657,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100111; Y = 7'b1010100; // Expected: {'Z': -1716}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100111; Y = 7'b1010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1658,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1716
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111010; Y = 7'b0110000; // Expected: {'Z': 2784}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111010; Y = 7'b0110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1659,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001010; Y = 7'b1100011; // Expected: {'Z': 1566}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001010; Y = 7'b1100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1660,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1566
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b1010111; // Expected: {'Z': 820}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b1010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1661,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000000; Y = 7'b1010110; // Expected: {'Z': 2688}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000000; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1662,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2688
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001000; Y = 7'b0100110; // Expected: {'Z': -2128}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001000; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1663,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000011; Y = 7'b0000011; // Expected: {'Z': -183}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000011; Y = 7'b0000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1664,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111001; Y = 7'b0000101; // Expected: {'Z': -35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111001; Y = 7'b0000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1665,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b0010111; // Expected: {'Z': -529}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b0010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1666,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -529
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001001; Y = 7'b1110000; // Expected: {'Z': 880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001001; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1667,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b0111101; // Expected: {'Z': -2074}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b0111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1668,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2074
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111110; Y = 7'b0001111; // Expected: {'Z': -30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111110; Y = 7'b0001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1669,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b1000011; // Expected: {'Z': -1037}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b1000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1670,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1037
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101010; Y = 7'b0100110; // Expected: {'Z': 1596}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101010; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1671,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1596
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001000; Y = 7'b0010000; // Expected: {'Z': -896}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001000; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1672,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110011; Y = 7'b1111010; // Expected: {'Z': 78}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110011; Y = 7'b1111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1673,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011111; Y = 7'b0000011; // Expected: {'Z': 93}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011111; Y = 7'b0000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1674,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000010; Y = 7'b0110110; // Expected: {'Z': 108}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000010; Y = 7'b0110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1675,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b1011110; // Expected: {'Z': -1802}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b1011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1676,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1802
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110000; Y = 7'b0000010; // Expected: {'Z': 96}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110000; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1677,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111100; Y = 7'b0000011; // Expected: {'Z': 180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111100; Y = 7'b0000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1678,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111001; Y = 7'b0110000; // Expected: {'Z': 2736}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111001; Y = 7'b0110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1679,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b0010011; // Expected: {'Z': -570}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b0010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1680,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -570
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001100; Y = 7'b0100010; // Expected: {'Z': -1768}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001100; Y = 7'b0100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1681,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1768
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010010; Y = 7'b0000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010010; Y = 7'b0000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1682,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101010; Y = 7'b0001101; // Expected: {'Z': -286}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101010; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1683,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -286
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b1010010; // Expected: {'Z': -46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b1010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1684,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001011; Y = 7'b1101001; // Expected: {'Z': 1219}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001011; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1685,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1219
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b1100110; // Expected: {'Z': -624}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b1100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1686,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b1000100; // Expected: {'Z': 2520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b1000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1687,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b0000101; // Expected: {'Z': -15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b0000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1688,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110000; Y = 7'b0001011; // Expected: {'Z': 528}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110000; Y = 7'b0001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1689,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001100; Y = 7'b0110101; // Expected: {'Z': -2756}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001100; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1690,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100111; Y = 7'b0100001; // Expected: {'Z': 1287}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100111; Y = 7'b0100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1691,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1287
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111010; Y = 7'b0000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111010; Y = 7'b0000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1692,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000010; Y = 7'b0011010; // Expected: {'Z': -1612}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000010; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1693,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110010; Y = 7'b1001000; // Expected: {'Z': 784}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110010; Y = 7'b1001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1694,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110011; Y = 7'b1010110; // Expected: {'Z': -2142}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110011; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1695,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011110; Y = 7'b1011100; // Expected: {'Z': -1080}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011110; Y = 7'b1011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1696,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100100; Y = 7'b0101001; // Expected: {'Z': 1476}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100100; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1697,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1476
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001011; Y = 7'b0011110; // Expected: {'Z': 330}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001011; Y = 7'b0011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1698,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 330
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100111; Y = 7'b1100010; // Expected: {'Z': 750}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100111; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1699,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b1100000; // Expected: {'Z': -1440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b1100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1700,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b1010000; // Expected: {'Z': 2016}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1701,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110101; Y = 7'b1000000; // Expected: {'Z': 704}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110101; Y = 7'b1000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1702,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 704
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b0101100; // Expected: {'Z': -660}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b0101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1703,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110110; Y = 7'b1101001; // Expected: {'Z': -1242}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110110; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1704,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b0000001; // Expected: {'Z': -30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b0000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1705,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111001; Y = 7'b1010101; // Expected: {'Z': 301}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111001; Y = 7'b1010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1706,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 301
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011001; Y = 7'b0001010; // Expected: {'Z': 250}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011001; Y = 7'b0001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1707,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111000; Y = 7'b1100010; // Expected: {'Z': -1680}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111000; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1708,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001110; Y = 7'b0110100; // Expected: {'Z': 728}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001110; Y = 7'b0110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1709,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100111; Y = 7'b1110110; // Expected: {'Z': 250}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100111; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1710,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b0101001; // Expected: {'Z': -1476}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1711,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1476
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b0011101; // Expected: {'Z': -1827}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1712,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1827
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b0101001; // Expected: {'Z': -697}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1713,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -697
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111100; Y = 7'b0110001; // Expected: {'Z': -196}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111100; Y = 7'b0110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1714,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110110; Y = 7'b0111010; // Expected: {'Z': 3132}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110110; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1715,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b0101100; // Expected: {'Z': -1012}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b0101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1716,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1012
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000111; Y = 7'b1110011; // Expected: {'Z': -91}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000111; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1717,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111001; Y = 7'b1010100; // Expected: {'Z': 308}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111001; Y = 7'b1010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1718,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 308
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100100; Y = 7'b1100100; // Expected: {'Z': -1008}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100100; Y = 7'b1100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1719,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b0011000; // Expected: {'Z': 72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b0011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1720,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010111; Y = 7'b0010001; // Expected: {'Z': -697}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010111; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1721,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -697
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b0010101; // Expected: {'Z': 1113}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b0010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1722,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001000; Y = 7'b0011001; // Expected: {'Z': -1400}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001000; Y = 7'b0011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1723,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010100; Y = 7'b0110101; // Expected: {'Z': -2332}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010100; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1724,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2332
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111000; Y = 7'b0010000; // Expected: {'Z': -128}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111000; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1725,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b1111000; // Expected: {'Z': -424}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b1111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1726,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -424
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101000; Y = 7'b0000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101000; Y = 7'b0000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1727,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b1010111; // Expected: {'Z': 1394}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b1010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1728,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1394
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110010; Y = 7'b0110011; // Expected: {'Z': 2550}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110010; Y = 7'b0110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1729,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110110; Y = 7'b0110100; // Expected: {'Z': 2808}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110110; Y = 7'b0110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1730,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b0011011; // Expected: {'Z': -972}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b0011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1731,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -972
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b0100110; // Expected: {'Z': -1292}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1732,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1292
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001110; Y = 7'b1100010; // Expected: {'Z': -420}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001110; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1733,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100010; Y = 7'b0100110; // Expected: {'Z': 1292}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100010; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1734,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1292
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100001; Y = 7'b1000010; // Expected: {'Z': 1922}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100001; Y = 7'b1000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1735,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1922
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b0101111; // Expected: {'Z': -1974}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b0101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1736,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1974
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110101; Y = 7'b0000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110101; Y = 7'b0000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1737,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b0001101; // Expected: {'Z': 221}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1738,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001100; Y = 7'b0100110; // Expected: {'Z': 456}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001100; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1739,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b0010011; // Expected: {'Z': 988}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b0010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1740,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 988
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b1100001; // Expected: {'Z': 1488}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b1100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1741,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101010; Y = 7'b1100010; // Expected: {'Z': -1260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101010; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1742,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b1101100; // Expected: {'Z': 800}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b1101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1743,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b0000110; // Expected: {'Z': -114}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b0000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1744,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101100; Y = 7'b0011100; // Expected: {'Z': 1232}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101100; Y = 7'b0011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1745,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b1111101; // Expected: {'Z': 54}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1746,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010011; Y = 7'b0001110; // Expected: {'Z': -630}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010011; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1747,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -630
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b1110010; // Expected: {'Z': 448}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b1110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1748,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 448
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110010; Y = 7'b1111010; // Expected: {'Z': 84}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110010; Y = 7'b1111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1749,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001100; Y = 7'b1111101; // Expected: {'Z': -36}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001100; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1750,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101011; Y = 7'b0110001; // Expected: {'Z': -1029}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101011; Y = 7'b0110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1751,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1029
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b0110001; // Expected: {'Z': -1568}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b0110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1752,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1568
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100101; Y = 7'b1101000; // Expected: {'Z': -888}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100101; Y = 7'b1101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1753,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111111; Y = 7'b0011010; // Expected: {'Z': 1638}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111111; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1754,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1638
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b1010110; // Expected: {'Z': 420}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1755,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110000; Y = 7'b1110010; // Expected: {'Z': 224}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110000; Y = 7'b1110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1756,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001011; Y = 7'b1100001; // Expected: {'Z': -341}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001011; Y = 7'b1100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1757,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -341
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010010; Y = 7'b0101100; // Expected: {'Z': 792}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010010; Y = 7'b0101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1758,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101011; Y = 7'b1111011; // Expected: {'Z': -215}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101011; Y = 7'b1111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1759,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -215
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b0000101; // Expected: {'Z': 120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b0000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1760,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b1011100; // Expected: {'Z': 648}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b1011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1761,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001001; Y = 7'b1111110; // Expected: {'Z': 110}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001001; Y = 7'b1111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1762,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b0100000; // Expected: {'Z': -896}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b0100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1763,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b0001100; // Expected: {'Z': -576}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b0001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1764,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101000; Y = 7'b1110100; // Expected: {'Z': 288}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101000; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1765,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001000; Y = 7'b0001000; // Expected: {'Z': -448}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001000; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1766,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -448
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b0000011; // Expected: {'Z': -120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b0000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1767,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b1110001; // Expected: {'Z': -675}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b1110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1768,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -675
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111000; Y = 7'b0111101; // Expected: {'Z': 3416}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111000; Y = 7'b0111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1769,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001110; Y = 7'b1111100; // Expected: {'Z': -56}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001110; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1770,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000011; Y = 7'b0001011; // Expected: {'Z': -671}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000011; Y = 7'b0001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1771,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -671
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111001; Y = 7'b0100000; // Expected: {'Z': 1824}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111001; Y = 7'b0100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1772,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1824
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b0110000; // Expected: {'Z': 144}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b0110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1773,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110111; Y = 7'b1100110; // Expected: {'Z': -1430}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110111; Y = 7'b1100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1774,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000100; Y = 7'b0101001; // Expected: {'Z': -2460}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000100; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1775,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2460
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b1110101; // Expected: {'Z': 330}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b1110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1776,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 330
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110001; Y = 7'b0100001; // Expected: {'Z': 1617}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110001; Y = 7'b0100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1777,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1617
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010010; Y = 7'b1111000; // Expected: {'Z': -144}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010010; Y = 7'b1111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1778,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011101; Y = 7'b0110001; // Expected: {'Z': -1715}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011101; Y = 7'b0110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1779,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1715
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b1001010; // Expected: {'Z': 540}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1780,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011101; Y = 7'b1011011; // Expected: {'Z': 1295}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011101; Y = 7'b1011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1781,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1295
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b1010111; // Expected: {'Z': 1394}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b1010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1782,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1394
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b0010001; // Expected: {'Z': -510}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1783,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -510
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b1110011; // Expected: {'Z': 442}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1784,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 442
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b0101110; // Expected: {'Z': -874}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b0101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1785,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -874
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000101; Y = 7'b0100010; // Expected: {'Z': -2006}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000101; Y = 7'b0100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1786,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2006
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b1101001; // Expected: {'Z': 345}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1787,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 345
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b1101101; // Expected: {'Z': -988}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b1101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1788,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -988
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101100; Y = 7'b0100000; // Expected: {'Z': 1408}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101100; Y = 7'b0100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1789,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101111; Y = 7'b0110111; // Expected: {'Z': 2585}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101111; Y = 7'b0110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1790,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2585
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111110; Y = 7'b1011010; // Expected: {'Z': 76}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111110; Y = 7'b1011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1791,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b0100000; // Expected: {'Z': 96}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b0100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1792,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011010; Y = 7'b1000000; // Expected: {'Z': -1664}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011010; Y = 7'b1000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1793,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1664
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b0011010; // Expected: {'Z': -1638}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1794,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1638
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b0111110; // Expected: {'Z': -62}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b0111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1795,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000000; Y = 7'b0011101; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000000; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1796,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b0001100; // Expected: {'Z': 636}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b0001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1797,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 636
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b0001010; // Expected: {'Z': -630}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b0001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1798,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -630
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b1010010; // Expected: {'Z': 1656}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b1010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1799,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1656
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010011; Y = 7'b1001110; // Expected: {'Z': -950}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010011; Y = 7'b1001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1800,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b0100000; // Expected: {'Z': 288}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b0100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1801,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010011; Y = 7'b0010001; // Expected: {'Z': 323}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010011; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1802,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 323
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110000; Y = 7'b1110111; // Expected: {'Z': -432}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110000; Y = 7'b1110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1803,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000011; Y = 7'b0101000; // Expected: {'Z': -2440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000011; Y = 7'b0101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1804,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011111; Y = 7'b0010010; // Expected: {'Z': 558}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011111; Y = 7'b0010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1805,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 558
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b1100101; // Expected: {'Z': -567}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1806,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -567
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010111; Y = 7'b1100101; // Expected: {'Z': -621}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010111; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1807,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -621
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101011; Y = 7'b0010000; // Expected: {'Z': 688}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101011; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1808,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 688
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100001; Y = 7'b1100011; // Expected: {'Z': 899}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100001; Y = 7'b1100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1809,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 899
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000011; Y = 7'b1100101; // Expected: {'Z': 1647}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000011; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1810,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1647
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b0001100; // Expected: {'Z': -180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b0001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1811,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b0010100; // Expected: {'Z': 180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b0010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1812,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b1010001; // Expected: {'Z': 1880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1813,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b0000010; // Expected: {'Z': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1814,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111001; Y = 7'b1111111; // Expected: {'Z': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111001; Y = 7'b1111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1815,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100000; Y = 7'b0001110; // Expected: {'Z': 448}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100000; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1816,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 448
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000110; Y = 7'b1110101; // Expected: {'Z': -66}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000110; Y = 7'b1110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1817,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011001; Y = 7'b1000110; // Expected: {'Z': -1450}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011001; Y = 7'b1000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1818,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101100; Y = 7'b1101110; // Expected: {'Z': -792}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101100; Y = 7'b1101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1819,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b1010110; // Expected: {'Z': 2016}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1820,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100101; Y = 7'b1100001; // Expected: {'Z': 837}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100101; Y = 7'b1100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1821,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 837
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001000; Y = 7'b1000111; // Expected: {'Z': -456}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001000; Y = 7'b1000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1822,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111010; Y = 7'b1010110; // Expected: {'Z': 252}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111010; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1823,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001101; Y = 7'b1100010; // Expected: {'Z': 1530}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001101; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1824,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1530
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010011; Y = 7'b1111111; // Expected: {'Z': 45}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010011; Y = 7'b1111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1825,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000111; Y = 7'b1000111; // Expected: {'Z': -399}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000111; Y = 7'b1000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1826,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -399
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010100; Y = 7'b0101101; // Expected: {'Z': -1980}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010100; Y = 7'b0101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1827,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010011; Y = 7'b1111010; // Expected: {'Z': -114}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010011; Y = 7'b1111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1828,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100010; Y = 7'b1101010; // Expected: {'Z': -748}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100010; Y = 7'b1101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1829,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -748
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110010; Y = 7'b1000100; // Expected: {'Z': -3000}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110010; Y = 7'b1000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1830,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101011; Y = 7'b1111001; // Expected: {'Z': 147}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101011; Y = 7'b1111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1831,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111011; Y = 7'b0010001; // Expected: {'Z': -85}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111011; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1832,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -85
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111011; Y = 7'b0010001; // Expected: {'Z': -85}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111011; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1833,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -85
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111001; Y = 7'b1000111; // Expected: {'Z': -3249}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111001; Y = 7'b1000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1834,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b0100111; // Expected: {'Z': -1404}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b0100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1835,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1404
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111010; Y = 7'b1011000; // Expected: {'Z': -2320}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111010; Y = 7'b1011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1836,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010010; Y = 7'b1010011; // Expected: {'Z': -810}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010010; Y = 7'b1010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1837,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -810
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001010; Y = 7'b1001111; // Expected: {'Z': -490}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001010; Y = 7'b1001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1838,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -490
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b1101100; // Expected: {'Z': -480}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b1101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1839,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010100; Y = 7'b1011010; // Expected: {'Z': 1672}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010100; Y = 7'b1011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1840,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010101; Y = 7'b0111000; // Expected: {'Z': -2408}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010101; Y = 7'b0111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1841,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001110; Y = 7'b1011111; // Expected: {'Z': -462}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001110; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1842,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b1111011; // Expected: {'Z': 180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b1111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1843,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000100; Y = 7'b0100111; // Expected: {'Z': 156}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000100; Y = 7'b0100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1844,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110011; Y = 7'b1110111; // Expected: {'Z': 117}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110011; Y = 7'b1110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1845,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001101; Y = 7'b0011010; // Expected: {'Z': -1326}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001101; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1846,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1326
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b1010001; // Expected: {'Z': -940}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1847,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -940
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111000; Y = 7'b1110100; // Expected: {'Z': 96}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111000; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1848,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001000; Y = 7'b0111100; // Expected: {'Z': 480}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001000; Y = 7'b0111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1849,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101011; Y = 7'b1101010; // Expected: {'Z': -946}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101011; Y = 7'b1101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1850,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -946
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110011; Y = 7'b1000101; // Expected: {'Z': -3009}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110011; Y = 7'b1000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1851,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3009
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b0000011; // Expected: {'Z': 72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b0000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1852,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111010; Y = 7'b1100010; // Expected: {'Z': 180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111010; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1853,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001100; Y = 7'b0111111; // Expected: {'Z': 756}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001100; Y = 7'b0111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1854,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010010; Y = 7'b1000100; // Expected: {'Z': 2760}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010010; Y = 7'b1000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1855,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b0001011; // Expected: {'Z': -187}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b0001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1856,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000000; Y = 7'b1110001; // Expected: {'Z': 960}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000000; Y = 7'b1110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1857,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101010; Y = 7'b1010100; // Expected: {'Z': -1848}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101010; Y = 7'b1010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1858,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b1101000; // Expected: {'Z': -408}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b1101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1859,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000101; Y = 7'b0111101; // Expected: {'Z': 305}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000101; Y = 7'b0111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1860,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 305
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010011; Y = 7'b1110010; // Expected: {'Z': -266}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010011; Y = 7'b1110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1861,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -266
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011110; Y = 7'b0010110; // Expected: {'Z': 660}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011110; Y = 7'b0010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1862,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001010; Y = 7'b0111011; // Expected: {'Z': 590}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001010; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1863,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 590
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011001; Y = 7'b1000010; // Expected: {'Z': 2418}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011001; Y = 7'b1000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1864,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2418
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100111; Y = 7'b0110111; // Expected: {'Z': -1375}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100111; Y = 7'b0110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1865,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1375
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b0100110; // Expected: {'Z': 1976}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1866,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1976
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111110; Y = 7'b0001001; // Expected: {'Z': -18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111110; Y = 7'b0001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1867,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b0010111; // Expected: {'Z': -69}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b0010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1868,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110101; Y = 7'b1010100; // Expected: {'Z': 484}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110101; Y = 7'b1010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1869,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 484
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110000; Y = 7'b1000111; // Expected: {'Z': -2736}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110000; Y = 7'b1000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1870,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b1100000; // Expected: {'Z': -544}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b1100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1871,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -544
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b0101110; // Expected: {'Z': -1932}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b0101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1872,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1932
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110011; Y = 7'b1100101; // Expected: {'Z': 351}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110011; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1873,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 351
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001111; Y = 7'b1111111; // Expected: {'Z': -15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001111; Y = 7'b1111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1874,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b1110000; // Expected: {'Z': 768}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1875,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 768
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b1011111; // Expected: {'Z': 1584}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1876,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1584
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001011; Y = 7'b0100110; // Expected: {'Z': 418}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001011; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1877,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 418
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100011; Y = 7'b1000001; // Expected: {'Z': 1827}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100011; Y = 7'b1000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1878,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1827
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b1100010; // Expected: {'Z': -720}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1879,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001000; Y = 7'b0000001; // Expected: {'Z': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001000; Y = 7'b0000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1880,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111100; Y = 7'b0000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111100; Y = 7'b0000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1881,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010110; Y = 7'b0000001; // Expected: {'Z': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010110; Y = 7'b0000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1882,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011001; Y = 7'b0000100; // Expected: {'Z': -156}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011001; Y = 7'b0000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1883,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011001; Y = 7'b1110001; // Expected: {'Z': -375}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011001; Y = 7'b1110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1884,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -375
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000110; Y = 7'b1111001; // Expected: {'Z': -42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000110; Y = 7'b1111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1885,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011111; Y = 7'b0010100; // Expected: {'Z': 620}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011111; Y = 7'b0010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1886,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111001; Y = 7'b1011100; // Expected: {'Z': -2052}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111001; Y = 7'b1011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1887,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2052
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100110; Y = 7'b0111111; // Expected: {'Z': -1638}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100110; Y = 7'b0111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1888,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1638
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111100; Y = 7'b0111001; // Expected: {'Z': -228}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111100; Y = 7'b0111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1889,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b0000110; // Expected: {'Z': 126}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b0000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1890,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b1111101; // Expected: {'Z': 126}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1891,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000111; Y = 7'b0111011; // Expected: {'Z': -3363}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000111; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1892,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3363
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100100; Y = 7'b0101111; // Expected: {'Z': 1692}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100100; Y = 7'b0101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1893,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1692
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b0100010; // Expected: {'Z': -1088}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b0100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1894,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1088
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101010; Y = 7'b1101110; // Expected: {'Z': -756}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101010; Y = 7'b1101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1895,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001010; Y = 7'b0101001; // Expected: {'Z': -2214}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001010; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1896,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101011; Y = 7'b1010100; // Expected: {'Z': -1892}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101011; Y = 7'b1010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1897,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1892
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111100; Y = 7'b0101000; // Expected: {'Z': -160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111100; Y = 7'b0101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1898,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011100; Y = 7'b1001101; // Expected: {'Z': -1428}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011100; Y = 7'b1001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1899,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1428
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000000; Y = 7'b1101110; // Expected: {'Z': 1152}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000000; Y = 7'b1101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1900,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001010; Y = 7'b0011111; // Expected: {'Z': -1674}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001010; Y = 7'b0011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1901,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1674
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011001; Y = 7'b0100010; // Expected: {'Z': 850}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011001; Y = 7'b0100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1902,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 850
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011110; Y = 7'b1101100; // Expected: {'Z': -600}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011110; Y = 7'b1101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1903,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b1000011; // Expected: {'Z': -2745}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b1000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1904,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2745
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110101; Y = 7'b1110000; // Expected: {'Z': 176}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110101; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1905,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010111; Y = 7'b1001110; // Expected: {'Z': -1150}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010111; Y = 7'b1001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1906,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b1111001; // Expected: {'Z': 224}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b1111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1907,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b0000011; // Expected: {'Z': 63}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b0000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1908,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b0001111; // Expected: {'Z': -270}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b0001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1909,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -270
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b1100010; // Expected: {'Z': -510}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1910,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -510
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b1001100; // Expected: {'Z': 1040}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b1001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1911,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b0000110; // Expected: {'Z': -192}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b0000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1912,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b0100100; // Expected: {'Z': -648}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b0100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1913,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b1100010; // Expected: {'Z': 300}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1914,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001010; Y = 7'b1010001; // Expected: {'Z': 2538}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001010; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1915,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2538
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010011; Y = 7'b0111010; // Expected: {'Z': -2610}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010011; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1916,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2610
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b0101000; // Expected: {'Z': 800}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b0101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1917,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011110; Y = 7'b0111010; // Expected: {'Z': 1740}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011110; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1918,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1740
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110001; Y = 7'b0011010; // Expected: {'Z': 1274}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110001; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1919,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1274
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000100; Y = 7'b1010101; // Expected: {'Z': 2580}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000100; Y = 7'b1010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1920,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100001; Y = 7'b1011110; // Expected: {'Z': 1054}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100001; Y = 7'b1011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1921,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1054
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b0100100; // Expected: {'Z': -1728}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b0100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1922,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b1111100; // Expected: {'Z': -4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1923,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101010; Y = 7'b1110011; // Expected: {'Z': -546}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101010; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1924,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b0100011; // Expected: {'Z': -1260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b0100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1925,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001100; Y = 7'b0010100; // Expected: {'Z': 240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001100; Y = 7'b0010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1926,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101111; Y = 7'b1110110; // Expected: {'Z': -470}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101111; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1927,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -470
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110101; Y = 7'b1100111; // Expected: {'Z': 275}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110101; Y = 7'b1100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1928,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 275
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011111; Y = 7'b0000110; // Expected: {'Z': 186}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011111; Y = 7'b0000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1929,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111011; Y = 7'b1110010; // Expected: {'Z': 70}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111011; Y = 7'b1110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1930,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010101; Y = 7'b1000001; // Expected: {'Z': 2709}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010101; Y = 7'b1000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1931,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2709
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101000; Y = 7'b0001010; // Expected: {'Z': -240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101000; Y = 7'b0001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1932,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b1110111; // Expected: {'Z': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b1110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1933,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b1011000; // Expected: {'Z': -40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b1011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1934,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100110; Y = 7'b0111110; // Expected: {'Z': -1612}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100110; Y = 7'b0111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1935,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b1110100; // Expected: {'Z': 216}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1936,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b1111110; // Expected: {'Z': -42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b1111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1937,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111111; Y = 7'b1000011; // Expected: {'Z': -3843}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111111; Y = 7'b1000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1938,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3843
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001101; Y = 7'b1110101; // Expected: {'Z': 561}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001101; Y = 7'b1110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1939,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 561
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011111; Y = 7'b1111011; // Expected: {'Z': -155}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011111; Y = 7'b1111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1940,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110011; Y = 7'b0001111; // Expected: {'Z': -195}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110011; Y = 7'b0001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1941,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110110; Y = 7'b0111000; // Expected: {'Z': 3024}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110110; Y = 7'b0111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1942,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101011; Y = 7'b0100101; // Expected: {'Z': 1591}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101011; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1943,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1591
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100000; Y = 7'b1111101; // Expected: {'Z': -96}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100000; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1944,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000000; Y = 7'b0111111; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000000; Y = 7'b0111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1945,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100101; Y = 7'b1010000; // Expected: {'Z': -1776}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100101; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1946,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1776
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101010; Y = 7'b0101011; // Expected: {'Z': 1806}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101010; Y = 7'b0101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1947,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1806
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000000; Y = 7'b0110101; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000000; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1948,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100110; Y = 7'b0101100; // Expected: {'Z': -1144}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100110; Y = 7'b0101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1949,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011100; Y = 7'b0010111; // Expected: {'Z': 644}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011100; Y = 7'b0010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1950,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 644
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b0110011; // Expected: {'Z': 459}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b0110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1951,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 459
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b0111111; // Expected: {'Z': -2142}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b0111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1952,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b0110111; // Expected: {'Z': 1320}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b0110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1953,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100000; Y = 7'b0110011; // Expected: {'Z': 1632}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100000; Y = 7'b0110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1954,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1632
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101000; Y = 7'b0101001; // Expected: {'Z': -984}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101000; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1955,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -984
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101111; Y = 7'b0000010; // Expected: {'Z': 94}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101111; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1956,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011110; Y = 7'b1111100; // Expected: {'Z': -120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011110; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1957,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001101; Y = 7'b1000111; // Expected: {'Z': -741}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001101; Y = 7'b1000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1958,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -741
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101000; Y = 7'b0000100; // Expected: {'Z': 160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101000; Y = 7'b0000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1959,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011001; Y = 7'b0000101; // Expected: {'Z': 125}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011001; Y = 7'b0000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1960,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b0011011; // Expected: {'Z': 81}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b0011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1961,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b0000111; // Expected: {'Z': -70}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b0000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1962,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011110; Y = 7'b0100001; // Expected: {'Z': 990}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011110; Y = 7'b0100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1963,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 990
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b1011000; // Expected: {'Z': -2480}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b1011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1964,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b1001110; // Expected: {'Z': 3150}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b1001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1965,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100000; Y = 7'b1110111; // Expected: {'Z': -288}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100000; Y = 7'b1110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1966,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010001; Y = 7'b1110110; // Expected: {'Z': 470}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010001; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1967,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 470
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b1011111; // Expected: {'Z': -1485}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1968,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1485
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110011; Y = 7'b0010100; // Expected: {'Z': -260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110011; Y = 7'b0010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1969,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101010; Y = 7'b0110111; // Expected: {'Z': -1210}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101010; Y = 7'b0110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1970,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110001; Y = 7'b0000010; // Expected: {'Z': 98}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110001; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1971,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001100; Y = 7'b1100001; // Expected: {'Z': 1612}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001100; Y = 7'b1100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1972,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101011; Y = 7'b0111010; // Expected: {'Z': -1218}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101011; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1973,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b1110100; // Expected: {'Z': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1974,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010101; Y = 7'b1001100; // Expected: {'Z': 2236}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010101; Y = 7'b1001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1975,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101100; Y = 7'b1001010; // Expected: {'Z': -2376}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101100; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1976,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2376
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001100; Y = 7'b1010010; // Expected: {'Z': -552}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001100; Y = 7'b1010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1977,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b0011110; // Expected: {'Z': 90}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b0011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1978,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011010; Y = 7'b0010101; // Expected: {'Z': 546}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011010; Y = 7'b0010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1979,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000101; Y = 7'b1111110; // Expected: {'Z': 118}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000101; Y = 7'b1111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1980,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b1000011; // Expected: {'Z': -1281}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b1000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1981,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1281
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b0011101; // Expected: {'Z': -870}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1982,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -870
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011100; Y = 7'b1000110; // Expected: {'Z': -1624}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011100; Y = 7'b1000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1983,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000010; Y = 7'b0010011; // Expected: {'Z': -1178}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000010; Y = 7'b0010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1984,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010011; Y = 7'b1010111; // Expected: {'Z': -779}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010011; Y = 7'b1010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1985,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -779
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b1000110; // Expected: {'Z': 2436}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b1000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1986,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2436
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011011; Y = 7'b0100100; // Expected: {'Z': 972}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011011; Y = 7'b0100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1987,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 972
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b0101010; // Expected: {'Z': -840}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b0101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1988,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000101; Y = 7'b0011011; // Expected: {'Z': -1593}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000101; Y = 7'b0011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1989,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1593
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b0111010; // Expected: {'Z': 1218}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1990,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101001; Y = 7'b1010111; // Expected: {'Z': -1681}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101001; Y = 7'b1010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1991,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1681
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100101; Y = 7'b1110011; // Expected: {'Z': 351}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100101; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1992,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 351
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b1001001; // Expected: {'Z': 660}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b1001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1993,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100100; Y = 7'b1111000; // Expected: {'Z': -288}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100100; Y = 7'b1111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1994,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101110; Y = 7'b1101001; // Expected: {'Z': -1058}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101110; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1995,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1058
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010000; Y = 7'b1000100; // Expected: {'Z': -960}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010000; Y = 7'b1000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1996,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b1010110; // Expected: {'Z': 1176}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1997,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000111; Y = 7'b0000101; // Expected: {'Z': 35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000111; Y = 7'b0000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1998,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b1001111; // Expected: {'Z': 3087}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b1001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1999,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3087
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111111; Y = 7'b1101011; // Expected: {'Z': -1323}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111111; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2000,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1323
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b0000010; // Expected: {'Z': 106}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2001,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001011; Y = 7'b0100001; // Expected: {'Z': 363}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001011; Y = 7'b0100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2002,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 363
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b1010000; // Expected: {'Z': -1152}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2003,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b0110110; // Expected: {'Z': 1296}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b0110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2004,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b0110110; // Expected: {'Z': -3402}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b0110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2005,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3402
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000000; Y = 7'b1000000; // Expected: {'Z': 4096}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000000; Y = 7'b1000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2006,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4096
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b1000000; // Expected: {'Z': 1472}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b1000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2007,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1472
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110001; Y = 7'b1111111; // Expected: {'Z': -49}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110001; Y = 7'b1111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2008,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b1000101; // Expected: {'Z': 1888}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b1000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2009,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100110; Y = 7'b1001100; // Expected: {'Z': 1352}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100110; Y = 7'b1001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2010,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100001; Y = 7'b0100000; // Expected: {'Z': -992}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100001; Y = 7'b0100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2011,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -992
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001110; Y = 7'b1001110; // Expected: {'Z': 2500}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001110; Y = 7'b1001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2012,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b0010001; // Expected: {'Z': -170}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2013,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b1010000; // Expected: {'Z': -2976}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2014,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2976
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b0110000; // Expected: {'Z': -480}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b0110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2015,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001010; Y = 7'b0000111; // Expected: {'Z': 70}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001010; Y = 7'b0000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2016,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b1101001; // Expected: {'Z': -552}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2017,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b1000101; // Expected: {'Z': -177}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b1000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2018,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -177
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b1001110; // Expected: {'Z': -1200}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b1001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2019,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111100; Y = 7'b1011000; // Expected: {'Z': -2400}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111100; Y = 7'b1011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2020,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b1011111; // Expected: {'Z': 627}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2021,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 627
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101010; Y = 7'b1101110; // Expected: {'Z': -756}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101010; Y = 7'b1101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2022,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000111; Y = 7'b1001010; // Expected: {'Z': 3078}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000111; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2023,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3078
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100110; Y = 7'b0000011; // Expected: {'Z': 114}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100110; Y = 7'b0000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2024,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000000; Y = 7'b0001110; // Expected: {'Z': -896}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000000; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2025,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000111; Y = 7'b1110101; // Expected: {'Z': -77}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000111; Y = 7'b1110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2026,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -77
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b1010100; // Expected: {'Z': 440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b1010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2027,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101010; Y = 7'b1010001; // Expected: {'Z': 1034}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101010; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2028,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1034
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b1000010; // Expected: {'Z': 1426}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b1000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2029,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1426
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b0100001; // Expected: {'Z': 693}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b0100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2030,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 693
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b0111001; // Expected: {'Z': -1596}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b0111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2031,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1596
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b0011011; // Expected: {'Z': -756}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b0011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2032,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110001; Y = 7'b1111001; // Expected: {'Z': -343}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110001; Y = 7'b1111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2033,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -343
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001010; Y = 7'b1101110; // Expected: {'Z': 972}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001010; Y = 7'b1101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2034,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 972
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b1101111; // Expected: {'Z': 612}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b1101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2035,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b1000000; // Expected: {'Z': -64}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b1000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2036,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011111; Y = 7'b0100001; // Expected: {'Z': -1089}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011111; Y = 7'b0100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2037,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1089
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b1101101; // Expected: {'Z': -57}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b1101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2038,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110011; Y = 7'b0110000; // Expected: {'Z': 2448}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110011; Y = 7'b0110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2039,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2448
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010001; Y = 7'b1011110; // Expected: {'Z': 1598}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010001; Y = 7'b1011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2040,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1598
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011110; Y = 7'b0001000; // Expected: {'Z': 240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011110; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2041,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010010; Y = 7'b0110100; // Expected: {'Z': 936}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010010; Y = 7'b0110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2042,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 936
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110101; Y = 7'b0010110; // Expected: {'Z': -242}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110101; Y = 7'b0010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2043,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101000; Y = 7'b0011000; // Expected: {'Z': -576}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101000; Y = 7'b0011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2044,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b1011001; // Expected: {'Z': -780}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b1011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2045,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101001; Y = 7'b1100000; // Expected: {'Z': -1312}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101001; Y = 7'b1100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2046,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1312
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001011; Y = 7'b1100000; // Expected: {'Z': -352}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001011; Y = 7'b1100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2047,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b0100100; // Expected: {'Z': -2268}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b0100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2048,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2268
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001001; Y = 7'b1111010; // Expected: {'Z': 330}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001001; Y = 7'b1111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2049,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 330
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001010; Y = 7'b1110000; // Expected: {'Z': -160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001010; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2050,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000000; Y = 7'b0000010; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000000; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2051,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000000; Y = 7'b0001001; // Expected: {'Z': -576}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000000; Y = 7'b0001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2052,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010101; Y = 7'b0111101; // Expected: {'Z': -2623}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010101; Y = 7'b0111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2053,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2623
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b0001010; // Expected: {'Z': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b0001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2054,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b0110111; // Expected: {'Z': 1100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b0110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2055,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001000; Y = 7'b0101100; // Expected: {'Z': -2464}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001000; Y = 7'b0101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2056,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011010; Y = 7'b0100001; // Expected: {'Z': 858}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011010; Y = 7'b0100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2057,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 858
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b0101000; // Expected: {'Z': -600}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b0101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2058,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000000; Y = 7'b0000100; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000000; Y = 7'b0000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2059,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110000; Y = 7'b0110011; // Expected: {'Z': -816}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110000; Y = 7'b0110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2060,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000010; Y = 7'b1010110; // Expected: {'Z': -84}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000010; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2061,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b0110101; // Expected: {'Z': -530}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2062,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -530
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000000; Y = 7'b1000101; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000000; Y = 7'b1000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2063,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b1111110; // Expected: {'Z': -2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b1111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2064,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100011; Y = 7'b1110001; // Expected: {'Z': 435}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100011; Y = 7'b1110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2065,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 435
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111101; Y = 7'b1010110; // Expected: {'Z': -2562}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111101; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2066,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2562
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b1011111; // Expected: {'Z': 924}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2067,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 924
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001000; Y = 7'b1010011; // Expected: {'Z': 2520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001000; Y = 7'b1010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2068,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010000; Y = 7'b1100001; // Expected: {'Z': -496}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010000; Y = 7'b1100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2069,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101000; Y = 7'b1110111; // Expected: {'Z': -360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101000; Y = 7'b1110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2070,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b1010001; // Expected: {'Z': 2961}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2071,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2961
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b0011111; // Expected: {'Z': -372}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b0011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2072,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -372
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b0011000; // Expected: {'Z': -816}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b0011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2073,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b0000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b0000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2074,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b0101011; // Expected: {'Z': -430}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b0101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2075,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100110; Y = 7'b1010101; // Expected: {'Z': 1118}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100110; Y = 7'b1010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2076,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b1000011; // Expected: {'Z': 1403}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b1000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2077,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1403
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110000; Y = 7'b0001011; // Expected: {'Z': 528}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110000; Y = 7'b0001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2078,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100000; Y = 7'b0101111; // Expected: {'Z': 1504}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100000; Y = 7'b0101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2079,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b0101110; // Expected: {'Z': -46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b0101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2080,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b0100010; // Expected: {'Z': -102}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b0100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2081,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b0100001; // Expected: {'Z': -1188}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b0100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2082,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100111; Y = 7'b0100110; // Expected: {'Z': -950}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100111; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2083,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100011; Y = 7'b1011010; // Expected: {'Z': 1102}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100011; Y = 7'b1011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2084,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100001; Y = 7'b1000100; // Expected: {'Z': 1860}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100001; Y = 7'b1000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2085,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1860
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010111; Y = 7'b1100111; // Expected: {'Z': -575}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010111; Y = 7'b1100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2086,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -575
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001000; Y = 7'b1011110; // Expected: {'Z': -272}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001000; Y = 7'b1011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2087,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -272
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b0010001; // Expected: {'Z': 884}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2088,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 884
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111011; Y = 7'b1010010; // Expected: {'Z': -2714}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111011; Y = 7'b1010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2089,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2714
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111011; Y = 7'b1100001; // Expected: {'Z': -1829}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111011; Y = 7'b1100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2090,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1829
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000101; Y = 7'b1001100; // Expected: {'Z': -260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000101; Y = 7'b1001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2091,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100110; Y = 7'b1011000; // Expected: {'Z': 1040}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100110; Y = 7'b1011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2092,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100101; Y = 7'b1111001; // Expected: {'Z': -259}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100101; Y = 7'b1111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2093,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -259
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101001; Y = 7'b1011001; // Expected: {'Z': -1599}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101001; Y = 7'b1011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2094,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1599
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001000; Y = 7'b1010100; // Expected: {'Z': 2464}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001000; Y = 7'b1010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2095,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011010; Y = 7'b1000010; // Expected: {'Z': 2356}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011010; Y = 7'b1000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2096,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2356
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000010; Y = 7'b1111001; // Expected: {'Z': -14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000010; Y = 7'b1111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2097,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111011; Y = 7'b1110111; // Expected: {'Z': -531}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111011; Y = 7'b1110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2098,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -531
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110101; Y = 7'b0110010; // Expected: {'Z': -550}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110101; Y = 7'b0110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2099,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001011; Y = 7'b1001010; // Expected: {'Z': -594}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001011; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2100,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -594
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b1100111; // Expected: {'Z': -500}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b1100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2101,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111000; Y = 7'b1111010; // Expected: {'Z': -336}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111000; Y = 7'b1111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2102,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -336
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011010; Y = 7'b0000100; // Expected: {'Z': 104}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011010; Y = 7'b0000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2103,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001001; Y = 7'b0111010; // Expected: {'Z': -3190}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001001; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2104,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000100; Y = 7'b1010000; // Expected: {'Z': 2880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000100; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2105,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010100; Y = 7'b0101110; // Expected: {'Z': -2024}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010100; Y = 7'b0101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2106,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011101; Y = 7'b1101111; // Expected: {'Z': 595}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011101; Y = 7'b1101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2107,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 595
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010010; Y = 7'b0001101; // Expected: {'Z': -598}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010010; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2108,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -598
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b1011000; // Expected: {'Z': 2520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b1011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2109,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001110; Y = 7'b1010110; // Expected: {'Z': 2100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001110; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2110,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111110; Y = 7'b0010001; // Expected: {'Z': -34}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111110; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2111,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011111; Y = 7'b1110101; // Expected: {'Z': -341}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011111; Y = 7'b1110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2112,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -341
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b1111100; // Expected: {'Z': -4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2113,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001011; Y = 7'b0010010; // Expected: {'Z': 198}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001011; Y = 7'b0010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2114,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101011; Y = 7'b0000010; // Expected: {'Z': -42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101011; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2115,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010100; Y = 7'b0001001; // Expected: {'Z': -396}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010100; Y = 7'b0001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2116,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -396
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100011; Y = 7'b1010011; // Expected: {'Z': 1305}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100011; Y = 7'b1010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2117,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1305
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000101; Y = 7'b1001010; // Expected: {'Z': 3186}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000101; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2118,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010011; Y = 7'b0100100; // Expected: {'Z': -1620}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010011; Y = 7'b0100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2119,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b0111011; // Expected: {'Z': -1357}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2120,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1357
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111000; Y = 7'b0001001; // Expected: {'Z': 504}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111000; Y = 7'b0001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2121,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b0100001; // Expected: {'Z': 1485}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b0100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2122,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1485
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000111; Y = 7'b0000110; // Expected: {'Z': -342}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000111; Y = 7'b0000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2123,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -342
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b1000001; // Expected: {'Z': -1260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b1000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2124,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000011; Y = 7'b1111110; // Expected: {'Z': 122}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000011; Y = 7'b1111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2125,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101111; Y = 7'b0010110; // Expected: {'Z': 1034}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101111; Y = 7'b0010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2126,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1034
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b1111110; // Expected: {'Z': 38}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b1111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2127,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b0111011; // Expected: {'Z': -1121}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2128,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b0110101; // Expected: {'Z': 1272}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2129,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1272
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000011; Y = 7'b0100101; // Expected: {'Z': -2257}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000011; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2130,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2257
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111000; Y = 7'b1100100; // Expected: {'Z': 224}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111000; Y = 7'b1100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2131,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011111; Y = 7'b1000110; // Expected: {'Z': -1798}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011111; Y = 7'b1000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2132,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000110; Y = 7'b1011110; // Expected: {'Z': 1972}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000110; Y = 7'b1011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2133,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1972
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000000; Y = 7'b0100010; // Expected: {'Z': -2176}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000000; Y = 7'b0100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2134,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110000; Y = 7'b1010011; // Expected: {'Z': 720}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110000; Y = 7'b1010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2135,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110000; Y = 7'b0010001; // Expected: {'Z': 816}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110000; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2136,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001100; Y = 7'b1001010; // Expected: {'Z': -648}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001100; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2137,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111000; Y = 7'b1000100; // Expected: {'Z': -3360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111000; Y = 7'b1000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2138,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b1110011; // Expected: {'Z': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2139,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b0101110; // Expected: {'Z': 46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b0101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2140,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101000; Y = 7'b0011000; // Expected: {'Z': 960}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101000; Y = 7'b0011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2141,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111100; Y = 7'b0111001; // Expected: {'Z': -228}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111100; Y = 7'b0111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2142,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011011; Y = 7'b1101101; // Expected: {'Z': -513}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011011; Y = 7'b1101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2143,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -513
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b0101101; // Expected: {'Z': 45}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b0101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2144,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001110; Y = 7'b0100011; // Expected: {'Z': -1750}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001110; Y = 7'b0100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2145,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b1001011; // Expected: {'Z': 1802}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b1001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2146,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1802
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b0010000; // Expected: {'Z': 336}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2147,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 336
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111001; Y = 7'b1001010; // Expected: {'Z': 378}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111001; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2148,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 378
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110111; Y = 7'b1011111; // Expected: {'Z': 297}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110111; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2149,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 297
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011011; Y = 7'b0101010; // Expected: {'Z': 1134}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011011; Y = 7'b0101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2150,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111011; Y = 7'b0010101; // Expected: {'Z': 1239}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111011; Y = 7'b0010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2151,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1239
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b0011111; // Expected: {'Z': -589}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b0011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2152,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -589
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b0010001; // Expected: {'Z': 765}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2153,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 765
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110010; Y = 7'b0111010; // Expected: {'Z': 2900}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110010; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2154,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101010; Y = 7'b0100001; // Expected: {'Z': 1386}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101010; Y = 7'b0100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2155,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1386
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001001; Y = 7'b1100001; // Expected: {'Z': 1705}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001001; Y = 7'b1100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2156,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1705
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001011; Y = 7'b0100111; // Expected: {'Z': -2067}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001011; Y = 7'b0100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2157,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2067
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010111; Y = 7'b1000011; // Expected: {'Z': 2501}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010111; Y = 7'b1000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2158,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2501
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110000; Y = 7'b0001001; // Expected: {'Z': 432}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110000; Y = 7'b0001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2159,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b0000010; // Expected: {'Z': -84}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2160,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001011; Y = 7'b0110001; // Expected: {'Z': -2597}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001011; Y = 7'b0110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2161,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2597
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b1111101; // Expected: {'Z': 60}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2162,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b1101010; // Expected: {'Z': 330}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b1101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2163,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 330
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011010; Y = 7'b0110010; // Expected: {'Z': -1900}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011010; Y = 7'b0110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2164,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100001; Y = 7'b1111001; // Expected: {'Z': -231}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100001; Y = 7'b1111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2165,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001111; Y = 7'b0000010; // Expected: {'Z': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001111; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2166,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100001; Y = 7'b0111000; // Expected: {'Z': 1848}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100001; Y = 7'b0111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2167,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010010; Y = 7'b1001100; // Expected: {'Z': 2392}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010010; Y = 7'b1001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2168,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100010; Y = 7'b1100101; // Expected: {'Z': -918}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100010; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2169,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -918
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001011; Y = 7'b0001000; // Expected: {'Z': -424}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001011; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2170,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -424
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101000; Y = 7'b0011000; // Expected: {'Z': 960}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101000; Y = 7'b0011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2171,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111001; Y = 7'b0101111; // Expected: {'Z': 2679}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111001; Y = 7'b0101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2172,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2679
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b1001010; // Expected: {'Z': 1944}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2173,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b1110010; // Expected: {'Z': 882}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b1110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2174,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 882
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000101; Y = 7'b1001001; // Expected: {'Z': -275}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000101; Y = 7'b1001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2175,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -275
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011010; Y = 7'b1111101; // Expected: {'Z': -78}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011010; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2176,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b1110011; // Expected: {'Z': -585}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2177,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -585
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001000; Y = 7'b1010101; // Expected: {'Z': 2408}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001000; Y = 7'b1010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2178,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b0111101; // Expected: {'Z': -3843}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b0111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2179,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3843
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100101; Y = 7'b0111110; // Expected: {'Z': 2294}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100101; Y = 7'b0111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2180,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2294
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b0010000; // Expected: {'Z': -240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2181,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b0110110; // Expected: {'Z': 918}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b0110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2182,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 918
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001001; Y = 7'b1000000; // Expected: {'Z': 3520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001001; Y = 7'b1000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2183,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b1011111; // Expected: {'Z': 1386}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2184,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1386
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110000; Y = 7'b0001101; // Expected: {'Z': 624}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110000; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2185,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000111; Y = 7'b1100110; // Expected: {'Z': 1482}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000111; Y = 7'b1100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2186,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1482
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b0100011; // Expected: {'Z': -665}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b0100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2187,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -665
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110101; Y = 7'b0001111; // Expected: {'Z': -165}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110101; Y = 7'b0001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2188,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b1111011; // Expected: {'Z': 90}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b1111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2189,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010111; Y = 7'b0111101; // Expected: {'Z': -2501}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010111; Y = 7'b0111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2190,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2501
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110011; Y = 7'b0001000; // Expected: {'Z': 408}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110011; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2191,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001111; Y = 7'b1001010; // Expected: {'Z': 2646}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001111; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2192,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2646
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101100; Y = 7'b0010011; // Expected: {'Z': 836}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101100; Y = 7'b0010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2193,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 836
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100010; Y = 7'b1000110; // Expected: {'Z': -1972}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100010; Y = 7'b1000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2194,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1972
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011100; Y = 7'b0010100; // Expected: {'Z': 560}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011100; Y = 7'b0010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2195,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101011; Y = 7'b1111100; // Expected: {'Z': 84}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101011; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2196,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b0001101; // Expected: {'Z': -546}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2197,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001100; Y = 7'b1001100; // Expected: {'Z': -624}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001100; Y = 7'b1001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2198,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b0001000; // Expected: {'Z': -160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2199,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101010; Y = 7'b0000111; // Expected: {'Z': -154}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101010; Y = 7'b0000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2200,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b1001010; // Expected: {'Z': -2862}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2201,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2862
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011011; Y = 7'b1110011; // Expected: {'Z': -351}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011011; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2202,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -351
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111100; Y = 7'b0011010; // Expected: {'Z': -104}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111100; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2203,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010010; Y = 7'b0110011; // Expected: {'Z': -2346}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010010; Y = 7'b0110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2204,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2346
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011111; Y = 7'b1000101; // Expected: {'Z': -1829}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011111; Y = 7'b1000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2205,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1829
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011101; Y = 7'b0010111; // Expected: {'Z': -805}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011101; Y = 7'b0010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2206,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -805
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100110; Y = 7'b0101000; // Expected: {'Z': 1520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100110; Y = 7'b0101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2207,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001111; Y = 7'b0100110; // Expected: {'Z': 570}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001111; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2208,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 570
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100010; Y = 7'b0001111; // Expected: {'Z': 510}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100010; Y = 7'b0001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2209,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 510
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b1010100; // Expected: {'Z': -880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b1010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2210,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100011; Y = 7'b0110101; // Expected: {'Z': 1855}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100011; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2211,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1855
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101000; Y = 7'b0000001; // Expected: {'Z': 40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101000; Y = 7'b0000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2212,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110010; Y = 7'b0011010; // Expected: {'Z': -364}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110010; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2213,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100011; Y = 7'b0110000; // Expected: {'Z': 1680}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100011; Y = 7'b0110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2214,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001100; Y = 7'b1101001; // Expected: {'Z': 1196}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001100; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2215,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110010; Y = 7'b1000101; // Expected: {'Z': -2950}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110010; Y = 7'b1000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2216,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110010; Y = 7'b1111101; // Expected: {'Z': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110010; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2217,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011010; Y = 7'b1011010; // Expected: {'Z': 1444}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011010; Y = 7'b1011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2218,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1444
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111110; Y = 7'b0000100; // Expected: {'Z': -8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111110; Y = 7'b0000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2219,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b0110011; // Expected: {'Z': -867}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b0110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2220,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -867
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010100; Y = 7'b1100100; // Expected: {'Z': 1232}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010100; Y = 7'b1100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2221,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000110; Y = 7'b0100111; // Expected: {'Z': -2262}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000110; Y = 7'b0100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2222,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2262
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001100; Y = 7'b0101111; // Expected: {'Z': 564}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001100; Y = 7'b0101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2223,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 564
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111000; Y = 7'b0100001; // Expected: {'Z': 1848}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111000; Y = 7'b0100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2224,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110010; Y = 7'b1000011; // Expected: {'Z': -3050}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110010; Y = 7'b1000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2225,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100100; Y = 7'b1110010; // Expected: {'Z': -504}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100100; Y = 7'b1110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2226,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101111; Y = 7'b1000100; // Expected: {'Z': -2820}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101111; Y = 7'b1000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2227,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011010; Y = 7'b0101101; // Expected: {'Z': 1170}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011010; Y = 7'b0101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2228,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100110; Y = 7'b1001011; // Expected: {'Z': -2014}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100110; Y = 7'b1001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2229,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2014
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011001; Y = 7'b0001100; // Expected: {'Z': -468}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011001; Y = 7'b0001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2230,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -468
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010010; Y = 7'b0010100; // Expected: {'Z': -920}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010010; Y = 7'b0010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2231,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b1111101; // Expected: {'Z': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2232,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000111; Y = 7'b1101100; // Expected: {'Z': -140}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000111; Y = 7'b1101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2233,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b1110110; // Expected: {'Z': -530}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2234,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -530
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b1100000; // Expected: {'Z': 736}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b1100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2235,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001010; Y = 7'b0110101; // Expected: {'Z': -2862}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001010; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2236,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2862
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001000; Y = 7'b0011001; // Expected: {'Z': -1400}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001000; Y = 7'b0011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2237,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b1001010; // Expected: {'Z': -2808}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2238,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011110; Y = 7'b0100111; // Expected: {'Z': 1170}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011110; Y = 7'b0100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2239,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b0110110; // Expected: {'Z': -1728}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b0110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2240,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110000; Y = 7'b1010101; // Expected: {'Z': -2064}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110000; Y = 7'b1010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2241,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2064
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b1100110; // Expected: {'Z': -1612}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b1100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2242,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b1010110; // Expected: {'Z': -882}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2243,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -882
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011100; Y = 7'b0000001; // Expected: {'Z': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011100; Y = 7'b0000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2244,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b1001101; // Expected: {'Z': 1632}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b1001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2245,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1632
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b1000010; // Expected: {'Z': 2232}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b1000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2246,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011111; Y = 7'b1010111; // Expected: {'Z': 1353}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011111; Y = 7'b1010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2247,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1353
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001010; Y = 7'b1101000; // Expected: {'Z': 1296}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001010; Y = 7'b1101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2248,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000111; Y = 7'b1001111; // Expected: {'Z': -343}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000111; Y = 7'b1001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2249,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -343
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b1010101; // Expected: {'Z': -2279}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b1010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2250,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2279
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111011; Y = 7'b0101010; // Expected: {'Z': -210}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111011; Y = 7'b0101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2251,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111110; Y = 7'b0000101; // Expected: {'Z': -10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111110; Y = 7'b0000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2252,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111100; Y = 7'b0110010; // Expected: {'Z': 3000}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111100; Y = 7'b0110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2253,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111010; Y = 7'b1111101; // Expected: {'Z': -174}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111010; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2254,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110111; Y = 7'b0001110; // Expected: {'Z': 770}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110111; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2255,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 770
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b1100011; // Expected: {'Z': 87}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b1100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2256,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 87
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001011; Y = 7'b0011011; // Expected: {'Z': -1431}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001011; Y = 7'b0011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2257,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1431
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001001; Y = 7'b0000011; // Expected: {'Z': -165}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001001; Y = 7'b0000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2258,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000110; Y = 7'b0111011; // Expected: {'Z': -3422}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000110; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2259,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3422
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000111; Y = 7'b0001001; // Expected: {'Z': -513}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000111; Y = 7'b0001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2260,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -513
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100011; Y = 7'b0111100; // Expected: {'Z': -1740}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100011; Y = 7'b0111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2261,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1740
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110010; Y = 7'b1001010; // Expected: {'Z': -2700}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110010; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2262,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001111; Y = 7'b0000101; // Expected: {'Z': 75}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001111; Y = 7'b0000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2263,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001111; Y = 7'b0010010; // Expected: {'Z': -882}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001111; Y = 7'b0010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2264,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -882
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100001; Y = 7'b0111101; // Expected: {'Z': 2013}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100001; Y = 7'b0111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2265,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2013
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b0110101; // Expected: {'Z': -2120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2266,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011011; Y = 7'b1011111; // Expected: {'Z': -891}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011011; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2267,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -891
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110011; Y = 7'b0110110; // Expected: {'Z': 2754}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110011; Y = 7'b0110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2268,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2754
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b1010000; // Expected: {'Z': 960}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2269,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000010; Y = 7'b1000010; // Expected: {'Z': -124}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000010; Y = 7'b1000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2270,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b1011001; // Expected: {'Z': -936}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b1011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2271,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -936
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110110; Y = 7'b1011111; // Expected: {'Z': -1782}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110110; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2272,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1782
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011011; Y = 7'b0011010; // Expected: {'Z': -962}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011011; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2273,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -962
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110010; Y = 7'b0111000; // Expected: {'Z': 2800}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110010; Y = 7'b0111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2274,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000100; Y = 7'b1001111; // Expected: {'Z': -196}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000100; Y = 7'b1001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2275,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b0001010; // Expected: {'Z': -360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b0001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2276,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b1000010; // Expected: {'Z': 1426}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b1000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2277,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1426
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101011; Y = 7'b1110100; // Expected: {'Z': 252}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101011; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2278,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100110; Y = 7'b0100001; // Expected: {'Z': 1254}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100110; Y = 7'b0100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2279,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b0001111; // Expected: {'Z': 780}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b0001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2280,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001111; Y = 7'b1001000; // Expected: {'Z': -840}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001111; Y = 7'b1001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2281,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000000; Y = 7'b0011110; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000000; Y = 7'b0011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2282,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110110; Y = 7'b0010100; // Expected: {'Z': 1080}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110110; Y = 7'b0010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2283,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111110; Y = 7'b1111110; // Expected: {'Z': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111110; Y = 7'b1111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2284,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111010; Y = 7'b1001011; // Expected: {'Z': -3074}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111010; Y = 7'b1001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2285,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3074
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b0101011; // Expected: {'Z': -1720}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b0101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2286,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000100; Y = 7'b1011101; // Expected: {'Z': -140}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000100; Y = 7'b1011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2287,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b0100101; // Expected: {'Z': -555}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2288,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -555
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110001; Y = 7'b0111110; // Expected: {'Z': 3038}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110001; Y = 7'b0111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2289,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3038
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101001; Y = 7'b0101101; // Expected: {'Z': 1845}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101001; Y = 7'b0101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2290,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1845
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100101; Y = 7'b1111110; // Expected: {'Z': -74}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100101; Y = 7'b1111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2291,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001010; Y = 7'b0010010; // Expected: {'Z': -972}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001010; Y = 7'b0010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2292,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -972
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b1101000; // Expected: {'Z': -1248}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b1101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2293,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b1111011; // Expected: {'Z': -100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b1111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2294,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111011; Y = 7'b1000000; // Expected: {'Z': 320}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111011; Y = 7'b1000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2295,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100110; Y = 7'b0100110; // Expected: {'Z': 1444}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100110; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2296,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1444
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011001; Y = 7'b0001110; // Expected: {'Z': 350}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011001; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2297,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b1001000; // Expected: {'Z': -168}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b1001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2298,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010011; Y = 7'b1001010; // Expected: {'Z': -1026}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010011; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2299,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1026
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b0110001; // Expected: {'Z': 441}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b0110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2300,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 441
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001101; Y = 7'b1010000; // Expected: {'Z': -624}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001101; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2301,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010000; Y = 7'b1100011; // Expected: {'Z': -464}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010000; Y = 7'b1100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2302,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b0101001; // Expected: {'Z': -615}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2303,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -615
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b1101110; // Expected: {'Z': 360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b1101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2304,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000101; Y = 7'b1011110; // Expected: {'Z': -170}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000101; Y = 7'b1011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2305,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b1100110; // Expected: {'Z': 442}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b1100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2306,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 442
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110011; Y = 7'b0010001; // Expected: {'Z': 867}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110011; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2307,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 867
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b0000110; // Expected: {'Z': 372}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b0000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2308,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 372
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010010; Y = 7'b0000101; // Expected: {'Z': -230}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010010; Y = 7'b0000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2309,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001100; Y = 7'b1110010; // Expected: {'Z': 728}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001100; Y = 7'b1110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2310,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b0011011; // Expected: {'Z': -459}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b0011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2311,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -459
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b1001000; // Expected: {'Z': -3472}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b1001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2312,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3472
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000010; Y = 7'b0010001; // Expected: {'Z': 34}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000010; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2313,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b0001110; // Expected: {'Z': 336}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2314,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 336
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111100; Y = 7'b0000111; // Expected: {'Z': 420}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111100; Y = 7'b0000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2315,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011111; Y = 7'b0101110; // Expected: {'Z': 1426}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011111; Y = 7'b0101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2316,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1426
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101110; Y = 7'b0001111; // Expected: {'Z': 690}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101110; Y = 7'b0001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2317,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 690
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100010; Y = 7'b1010001; // Expected: {'Z': -1598}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100010; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2318,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1598
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010111; Y = 7'b0011111; // Expected: {'Z': -1271}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010111; Y = 7'b0011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2319,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1271
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b0000011; // Expected: {'Z': 159}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b0000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2320,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000101; Y = 7'b0100101; // Expected: {'Z': 185}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000101; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2321,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b1010101; // Expected: {'Z': -2236}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b1010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2322,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b0001001; // Expected: {'Z': -180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b0001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2323,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100011; Y = 7'b0010111; // Expected: {'Z': -667}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100011; Y = 7'b0010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2324,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -667
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110000; Y = 7'b0010100; // Expected: {'Z': -320}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110000; Y = 7'b0010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2325,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b1000101; // Expected: {'Z': 2360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b1000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2326,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000010; Y = 7'b1111010; // Expected: {'Z': -12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000010; Y = 7'b1111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2327,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111001; Y = 7'b1111100; // Expected: {'Z': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111001; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2328,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101011; Y = 7'b1001001; // Expected: {'Z': 1155}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101011; Y = 7'b1001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2329,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100101; Y = 7'b0100101; // Expected: {'Z': -999}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100101; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2330,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -999
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001010; Y = 7'b0101010; // Expected: {'Z': 420}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001010; Y = 7'b0101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2331,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111011; Y = 7'b0100111; // Expected: {'Z': -195}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111011; Y = 7'b0100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2332,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011110; Y = 7'b1010011; // Expected: {'Z': -1350}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011110; Y = 7'b1010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2333,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001110; Y = 7'b0000100; // Expected: {'Z': 56}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001110; Y = 7'b0000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2334,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011010; Y = 7'b1000101; // Expected: {'Z': -1534}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011010; Y = 7'b1000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2335,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1534
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110111; Y = 7'b0100101; // Expected: {'Z': -333}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110111; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2336,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -333
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110000; Y = 7'b1000001; // Expected: {'Z': 1008}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110000; Y = 7'b1000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2337,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001110; Y = 7'b1101111; // Expected: {'Z': -238}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001110; Y = 7'b1101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2338,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110111; Y = 7'b0010010; // Expected: {'Z': -162}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110111; Y = 7'b0010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2339,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111111; Y = 7'b1010111; // Expected: {'Z': -2583}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111111; Y = 7'b1010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2340,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2583
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100001; Y = 7'b0110101; // Expected: {'Z': 1749}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100001; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2341,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1749
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b1001011; // Expected: {'Z': 636}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b1001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2342,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 636
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100101; Y = 7'b0100011; // Expected: {'Z': -945}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100101; Y = 7'b0100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2343,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -945
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110010; Y = 7'b1000010; // Expected: {'Z': 868}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110010; Y = 7'b1000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2344,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 868
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001001; Y = 7'b1001011; // Expected: {'Z': 2915}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001001; Y = 7'b1001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2345,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2915
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001101; Y = 7'b1110000; // Expected: {'Z': -208}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001101; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2346,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011001; Y = 7'b1011110; // Expected: {'Z': -850}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011001; Y = 7'b1011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2347,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -850
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110011; Y = 7'b0010110; // Expected: {'Z': 1122}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110011; Y = 7'b0010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2348,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010000; Y = 7'b1100011; // Expected: {'Z': -464}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010000; Y = 7'b1100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2349,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b0101110; // Expected: {'Z': -690}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b0101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2350,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -690
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110011; Y = 7'b0110011; // Expected: {'Z': -663}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110011; Y = 7'b0110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2351,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -663
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001101; Y = 7'b0010000; // Expected: {'Z': 208}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001101; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2352,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100110; Y = 7'b1010001; // Expected: {'Z': 1222}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100110; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2353,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111000; Y = 7'b0001111; // Expected: {'Z': 840}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111000; Y = 7'b0001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2354,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110011; Y = 7'b0111111; // Expected: {'Z': -819}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110011; Y = 7'b0111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2355,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -819
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100110; Y = 7'b0000101; // Expected: {'Z': -130}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100110; Y = 7'b0000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2356,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111000; Y = 7'b0100101; // Expected: {'Z': -296}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111000; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2357,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b1100010; // Expected: {'Z': 1080}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2358,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101001; Y = 7'b0101100; // Expected: {'Z': 1804}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101001; Y = 7'b0101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2359,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1804
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011001; Y = 7'b0001010; // Expected: {'Z': 250}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011001; Y = 7'b0001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2360,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101000; Y = 7'b1101000; // Expected: {'Z': 576}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101000; Y = 7'b1101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2361,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100111; Y = 7'b1001111; // Expected: {'Z': 1225}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100111; Y = 7'b1001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2362,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100110; Y = 7'b1101011; // Expected: {'Z': -798}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100110; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2363,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101010; Y = 7'b1101001; // Expected: {'Z': 506}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101010; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2364,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 506
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111101; Y = 7'b0110111; // Expected: {'Z': 3355}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111101; Y = 7'b0110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2365,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3355
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111100; Y = 7'b0011001; // Expected: {'Z': -100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111100; Y = 7'b0011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2366,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010010; Y = 7'b1000111; // Expected: {'Z': 2622}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010010; Y = 7'b1000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2367,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2622
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110010; Y = 7'b0111110; // Expected: {'Z': 3100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110010; Y = 7'b0111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2368,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b0011101; // Expected: {'Z': -1392}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2369,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101111; Y = 7'b1011000; // Expected: {'Z': -1880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101111; Y = 7'b1011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2370,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111101; Y = 7'b0010010; // Expected: {'Z': 1098}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111101; Y = 7'b0010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2371,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1098
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b0010000; // Expected: {'Z': -576}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2372,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b1111011; // Expected: {'Z': 90}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b1111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2373,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b0011000; // Expected: {'Z': -1152}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b0011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2374,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010110; Y = 7'b0100101; // Expected: {'Z': 814}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010110; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2375,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 814
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111000; Y = 7'b1101101; // Expected: {'Z': -1064}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111000; Y = 7'b1101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2376,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1064
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110010; Y = 7'b1111011; // Expected: {'Z': -250}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110010; Y = 7'b1111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2377,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b1001010; // Expected: {'Z': 1620}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2378,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010000; Y = 7'b1000111; // Expected: {'Z': -912}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010000; Y = 7'b1000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2379,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -912
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b0001101; // Expected: {'Z': -468}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2380,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -468
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111001; Y = 7'b1100010; // Expected: {'Z': 210}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111001; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2381,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011001; Y = 7'b0000001; // Expected: {'Z': -39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011001; Y = 7'b0000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2382,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010010; Y = 7'b0001011; // Expected: {'Z': -506}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010010; Y = 7'b0001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2383,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -506
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b1100111; // Expected: {'Z': -225}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b1100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2384,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000000; Y = 7'b0000011; // Expected: {'Z': -192}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000000; Y = 7'b0000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2385,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011101; Y = 7'b0110111; // Expected: {'Z': 1595}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011101; Y = 7'b0110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2386,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1595
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b0011000; // Expected: {'Z': -768}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b0011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2387,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -768
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b0101110; // Expected: {'Z': 414}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b0101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2388,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 414
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010001; Y = 7'b1000100; // Expected: {'Z': 2820}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010001; Y = 7'b1000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2389,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000111; Y = 7'b0110010; // Expected: {'Z': -2850}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000111; Y = 7'b0110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2390,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2850
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111011; Y = 7'b1011111; // Expected: {'Z': 165}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111011; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2391,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011110; Y = 7'b1010101; // Expected: {'Z': -1290}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011110; Y = 7'b1010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2392,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1290
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111010; Y = 7'b0010000; // Expected: {'Z': 928}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111010; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2393,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 928
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110010; Y = 7'b0111000; // Expected: {'Z': -784}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110010; Y = 7'b0111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2394,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100110; Y = 7'b0110111; // Expected: {'Z': -1430}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100110; Y = 7'b0110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2395,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b1100110; // Expected: {'Z': 936}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b1100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2396,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 936
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011011; Y = 7'b0110011; // Expected: {'Z': 1377}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011011; Y = 7'b0110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2397,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1377
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b0101101; // Expected: {'Z': -1620}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b0101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2398,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b1011010; // Expected: {'Z': 1824}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b1011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2399,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1824
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b1101010; // Expected: {'Z': 264}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b1101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2400,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b0101010; // Expected: {'Z': 714}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b0101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2401,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 714
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b1011000; // Expected: {'Z': 920}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b1011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2402,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b0000010; // Expected: {'Z': 104}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2403,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010111; Y = 7'b0111101; // Expected: {'Z': 1403}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010111; Y = 7'b0111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2404,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1403
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010011; Y = 7'b0001000; // Expected: {'Z': 152}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010011; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2405,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b0110000; // Expected: {'Z': -2016}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b0110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2406,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111001; Y = 7'b0010000; // Expected: {'Z': 912}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111001; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2407,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 912
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b1110010; // Expected: {'Z': 392}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b1110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2408,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b1011001; // Expected: {'Z': -780}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b1011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2409,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101001; Y = 7'b0101100; // Expected: {'Z': 1804}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101001; Y = 7'b0101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2410,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1804
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101100; Y = 7'b0100110; // Expected: {'Z': 1672}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101100; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2411,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001011; Y = 7'b1010111; // Expected: {'Z': -451}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001011; Y = 7'b1010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2412,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -451
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110111; Y = 7'b1101001; // Expected: {'Z': -1265}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110111; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2413,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1265
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b1110011; // Expected: {'Z': 260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2414,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001000; Y = 7'b0010101; // Expected: {'Z': 168}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001000; Y = 7'b0010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2415,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010100; Y = 7'b1000011; // Expected: {'Z': 2684}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010100; Y = 7'b1000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2416,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2684
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101001; Y = 7'b1110101; // Expected: {'Z': -451}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101001; Y = 7'b1110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2417,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -451
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000100; Y = 7'b1111010; // Expected: {'Z': -24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000100; Y = 7'b1111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2418,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b1111100; // Expected: {'Z': 40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2419,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100101; Y = 7'b0011111; // Expected: {'Z': -837}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100101; Y = 7'b0011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2420,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -837
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b0011101; // Expected: {'Z': 1537}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2421,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1537
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000100; Y = 7'b1110110; // Expected: {'Z': -40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000100; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2422,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110000; Y = 7'b0001111; // Expected: {'Z': 720}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110000; Y = 7'b0001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2423,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000101; Y = 7'b1001000; // Expected: {'Z': 3304}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000101; Y = 7'b1001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2424,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3304
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001010; Y = 7'b0111001; // Expected: {'Z': -3078}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001010; Y = 7'b0111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2425,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3078
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b0110100; // Expected: {'Z': -1456}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b0110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2426,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001010; Y = 7'b1101101; // Expected: {'Z': -190}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001010; Y = 7'b1101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2427,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011001; Y = 7'b0010000; // Expected: {'Z': 400}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011001; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2428,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100000; Y = 7'b0110000; // Expected: {'Z': 1536}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100000; Y = 7'b0110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2429,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1536
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101011; Y = 7'b0011010; // Expected: {'Z': -546}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101011; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2430,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001111; Y = 7'b1010011; // Expected: {'Z': 2205}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001111; Y = 7'b1010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2431,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b0110011; // Expected: {'Z': -153}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b0110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2432,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -153
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010010; Y = 7'b1111110; // Expected: {'Z': 92}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010010; Y = 7'b1111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2433,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000110; Y = 7'b0000100; // Expected: {'Z': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000110; Y = 7'b0000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2434,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b1001010; // Expected: {'Z': 1026}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2435,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1026
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010101; Y = 7'b0101101; // Expected: {'Z': -1935}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010101; Y = 7'b0101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2436,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1935
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b1001011; // Expected: {'Z': 1484}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b1001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2437,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1484
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001111; Y = 7'b1011011; // Expected: {'Z': -555}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001111; Y = 7'b1011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2438,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -555
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010111; Y = 7'b0010110; // Expected: {'Z': 506}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010111; Y = 7'b0010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2439,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 506
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001001; Y = 7'b1100111; // Expected: {'Z': 1375}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001001; Y = 7'b1100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2440,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1375
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b1001111; // Expected: {'Z': -49}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b1001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2441,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001111; Y = 7'b0001101; // Expected: {'Z': 195}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001111; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2442,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000101; Y = 7'b0110011; // Expected: {'Z': 255}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000101; Y = 7'b0110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2443,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110101; Y = 7'b1000011; // Expected: {'Z': 671}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110101; Y = 7'b1000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2444,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 671
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100001; Y = 7'b1011100; // Expected: {'Z': 1116}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100001; Y = 7'b1011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2445,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011001; Y = 7'b0101000; // Expected: {'Z': -1560}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011001; Y = 7'b0101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2446,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b1011010; // Expected: {'Z': -1710}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b1011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2447,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1710
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001101; Y = 7'b1001001; // Expected: {'Z': 2805}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001101; Y = 7'b1001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2448,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2805
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000110; Y = 7'b0111111; // Expected: {'Z': 378}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000110; Y = 7'b0111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2449,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 378
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110000; Y = 7'b1000000; // Expected: {'Z': 1024}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110000; Y = 7'b1000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2450,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b0001110; // Expected: {'Z': 280}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2451,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100011; Y = 7'b1001001; // Expected: {'Z': -1925}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100011; Y = 7'b1001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2452,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1925
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001110; Y = 7'b1001010; // Expected: {'Z': -756}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001110; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2453,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011111; Y = 7'b1100100; // Expected: {'Z': -868}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011111; Y = 7'b1100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2454,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -868
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100001; Y = 7'b0011101; // Expected: {'Z': 957}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100001; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2455,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 957
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001000; Y = 7'b0101100; // Expected: {'Z': 352}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001000; Y = 7'b0101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2456,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001111; Y = 7'b1011111; // Expected: {'Z': -495}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001111; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2457,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -495
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010001; Y = 7'b1100001; // Expected: {'Z': 1457}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010001; Y = 7'b1100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2458,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1457
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111010; Y = 7'b1111000; // Expected: {'Z': -464}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111010; Y = 7'b1111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2459,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b0101000; // Expected: {'Z': -800}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b0101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2460,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110011; Y = 7'b0100111; // Expected: {'Z': -507}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110011; Y = 7'b0100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2461,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -507
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101000; Y = 7'b1100100; // Expected: {'Z': -1120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101000; Y = 7'b1100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2462,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b1110100; // Expected: {'Z': -204}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2463,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100001; Y = 7'b1000010; // Expected: {'Z': 1922}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100001; Y = 7'b1000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2464,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1922
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010010; Y = 7'b1100111; // Expected: {'Z': -450}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010010; Y = 7'b1100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2465,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010111; Y = 7'b1001111; // Expected: {'Z': 2009}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010111; Y = 7'b1001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2466,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2009
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111101; Y = 7'b0000011; // Expected: {'Z': 183}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111101; Y = 7'b0000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2467,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011101; Y = 7'b0101101; // Expected: {'Z': 1305}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011101; Y = 7'b0101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2468,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1305
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110000; Y = 7'b1011011; // Expected: {'Z': 592}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110000; Y = 7'b1011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2469,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 592
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b1001101; // Expected: {'Z': 1530}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b1001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2470,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1530
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b0010111; // Expected: {'Z': 460}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b0010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2471,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 460
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001111; Y = 7'b1110000; // Expected: {'Z': -240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001111; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2472,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110011; Y = 7'b0101001; // Expected: {'Z': -533}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110011; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2473,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -533
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b1101111; // Expected: {'Z': 255}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b1101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2474,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001000; Y = 7'b1110011; // Expected: {'Z': -104}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001000; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2475,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001010; Y = 7'b1111101; // Expected: {'Z': 162}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001010; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2476,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111001; Y = 7'b0011000; // Expected: {'Z': 1368}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111001; Y = 7'b0011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2477,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010011; Y = 7'b0101010; // Expected: {'Z': 798}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010011; Y = 7'b0101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2478,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101001; Y = 7'b1101111; // Expected: {'Z': -697}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101001; Y = 7'b1101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2479,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -697
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b1111011; // Expected: {'Z': 100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b1111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2480,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b0110100; // Expected: {'Z': 52}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b0110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2481,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011111; Y = 7'b1000001; // Expected: {'Z': 2079}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011111; Y = 7'b1000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2482,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2079
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100111; Y = 7'b0001001; // Expected: {'Z': 351}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100111; Y = 7'b0001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2483,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 351
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110000; Y = 7'b0101000; // Expected: {'Z': 1920}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110000; Y = 7'b0101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2484,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101011; Y = 7'b0011110; // Expected: {'Z': 1290}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101011; Y = 7'b0011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2485,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1290
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010010; Y = 7'b0100010; // Expected: {'Z': 612}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010010; Y = 7'b0100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2486,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010101; Y = 7'b0100010; // Expected: {'Z': -1462}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010101; Y = 7'b0100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2487,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b0110011; // Expected: {'Z': -1428}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b0110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2488,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1428
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011111; Y = 7'b0110110; // Expected: {'Z': 1674}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011111; Y = 7'b0110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2489,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1674
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110010; Y = 7'b0111011; // Expected: {'Z': -826}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110010; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2490,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -826
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000100; Y = 7'b1100010; // Expected: {'Z': 1800}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000100; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2491,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111010; Y = 7'b0011011; // Expected: {'Z': -162}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111010; Y = 7'b0011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2492,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001110; Y = 7'b1010010; // Expected: {'Z': -644}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001110; Y = 7'b1010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2493,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -644
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111000; Y = 7'b0110101; // Expected: {'Z': -424}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111000; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2494,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -424
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b0111111; // Expected: {'Z': 3339}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b0111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2495,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3339
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111110; Y = 7'b1101111; // Expected: {'Z': 34}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111110; Y = 7'b1101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2496,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111111; Y = 7'b0010001; // Expected: {'Z': 1071}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111111; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2497,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1071
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011001; Y = 7'b0100001; // Expected: {'Z': -1287}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011001; Y = 7'b0100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2498,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1287
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b1001101; // Expected: {'Z': -2652}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b1001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2499,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2652
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011101; Y = 7'b0001111; // Expected: {'Z': 435}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011101; Y = 7'b0001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2500,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 435
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001110; Y = 7'b0110011; // Expected: {'Z': -2550}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001110; Y = 7'b0110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2501,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101001; Y = 7'b0000110; // Expected: {'Z': 246}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101001; Y = 7'b0000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2502,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100001; Y = 7'b1100101; // Expected: {'Z': 837}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100001; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2503,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 837
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110000; Y = 7'b1111111; // Expected: {'Z': -48}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110000; Y = 7'b1111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2504,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010010; Y = 7'b1101110; // Expected: {'Z': 828}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010010; Y = 7'b1101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2505,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101010; Y = 7'b0100111; // Expected: {'Z': 1638}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101010; Y = 7'b0100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2506,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1638
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001110; Y = 7'b1000011; // Expected: {'Z': -854}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001110; Y = 7'b1000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2507,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -854
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b1000000; // Expected: {'Z': -192}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b1000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2508,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011011; Y = 7'b1100100; // Expected: {'Z': 1036}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011011; Y = 7'b1100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2509,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1036
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b1001010; // Expected: {'Z': -486}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2510,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -486
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011010; Y = 7'b0100111; // Expected: {'Z': 1014}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011010; Y = 7'b0100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2511,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1014
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010110; Y = 7'b1110110; // Expected: {'Z': -220}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010110; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2512,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110110; Y = 7'b0110101; // Expected: {'Z': 2862}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110110; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2513,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2862
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010001; Y = 7'b1110011; // Expected: {'Z': 611}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010001; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2514,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 611
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111010; Y = 7'b0000100; // Expected: {'Z': -24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111010; Y = 7'b0000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2515,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b1110010; // Expected: {'Z': -294}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b1110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2516,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -294
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001010; Y = 7'b0011100; // Expected: {'Z': 280}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001010; Y = 7'b0011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2517,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010110; Y = 7'b1001000; // Expected: {'Z': -1232}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010110; Y = 7'b1001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2518,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b0011101; // Expected: {'Z': 261}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2519,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 261
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111000; Y = 7'b1100100; // Expected: {'Z': 224}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111000; Y = 7'b1100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2520,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001100; Y = 7'b0111110; // Expected: {'Z': -3224}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001100; Y = 7'b0111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2521,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b0011100; // Expected: {'Z': 672}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b0011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2522,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011110; Y = 7'b1000111; // Expected: {'Z': -1710}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011110; Y = 7'b1000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2523,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1710
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b0001010; // Expected: {'Z': 240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b0001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2524,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b0100110; // Expected: {'Z': -760}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2525,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101010; Y = 7'b0110110; // Expected: {'Z': 2268}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101010; Y = 7'b0110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2526,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2268
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101000; Y = 7'b0011011; // Expected: {'Z': -648}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101000; Y = 7'b0011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2527,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100011; Y = 7'b0101101; // Expected: {'Z': 1575}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100011; Y = 7'b0101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2528,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1575
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b1011101; // Expected: {'Z': 2205}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b1011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2529,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b0011111; // Expected: {'Z': -558}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b0011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2530,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -558
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111111; Y = 7'b0011110; // Expected: {'Z': 1890}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111111; Y = 7'b0011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2531,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1890
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001100; Y = 7'b0111100; // Expected: {'Z': 720}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001100; Y = 7'b0111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2532,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b0011101; // Expected: {'Z': -1827}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2533,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1827
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111001; Y = 7'b1011111; // Expected: {'Z': -1881}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111001; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2534,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1881
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001111; Y = 7'b0011010; // Expected: {'Z': -1274}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001111; Y = 7'b0011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2535,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1274
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001000; Y = 7'b0100010; // Expected: {'Z': -1904}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001000; Y = 7'b0100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2536,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1904
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b0011001; // Expected: {'Z': -300}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b0011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2537,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100110; Y = 7'b1010011; // Expected: {'Z': 1170}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100110; Y = 7'b1010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2538,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011111; Y = 7'b1001110; // Expected: {'Z': 1650}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011111; Y = 7'b1001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2539,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b1110000; // Expected: {'Z': -384}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2540,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -384
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b1010101; // Expected: {'Z': -731}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b1010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2541,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -731
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110011; Y = 7'b1100100; // Expected: {'Z': -1428}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110011; Y = 7'b1100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2542,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1428
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110110; Y = 7'b1011001; // Expected: {'Z': -2106}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110110; Y = 7'b1011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2543,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111001; Y = 7'b1011101; // Expected: {'Z': -1995}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111001; Y = 7'b1011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2544,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1995
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b1111111; // Expected: {'Z': -24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b1111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2545,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b0101011; // Expected: {'Z': 43}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b0101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2546,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010111; Y = 7'b0110111; // Expected: {'Z': -2255}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010111; Y = 7'b0110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2547,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100101; Y = 7'b0010011; // Expected: {'Z': -513}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100101; Y = 7'b0010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2548,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -513
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b1110001; // Expected: {'Z': 945}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b1110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2549,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 945
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011011; Y = 7'b1101101; // Expected: {'Z': -513}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011011; Y = 7'b1101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2550,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -513
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111001; Y = 7'b1011001; // Expected: {'Z': 273}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111001; Y = 7'b1011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2551,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 273
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110011; Y = 7'b0001101; // Expected: {'Z': 663}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110011; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2552,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 663
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b0101101; // Expected: {'Z': 2790}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b0101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2553,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2790
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000000; Y = 7'b0010101; // Expected: {'Z': -1344}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000000; Y = 7'b0010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2554,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1344
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101001; Y = 7'b0001100; // Expected: {'Z': 492}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101001; Y = 7'b0001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2555,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 492
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100111; Y = 7'b1011110; // Expected: {'Z': 850}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100111; Y = 7'b1011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2556,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 850
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001111; Y = 7'b0011110; // Expected: {'Z': 450}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001111; Y = 7'b0011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2557,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110000; Y = 7'b1000000; // Expected: {'Z': -3072}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110000; Y = 7'b1000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2558,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3072
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101000; Y = 7'b1010000; // Expected: {'Z': 1152}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101000; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2559,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001110; Y = 7'b0001110; // Expected: {'Z': 196}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001110; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2560,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001111; Y = 7'b1110001; // Expected: {'Z': -225}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001111; Y = 7'b1110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2561,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b1111111; // Expected: {'Z': 40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b1111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2562,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b0100010; // Expected: {'Z': -1088}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b0100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2563,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1088
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011010; Y = 7'b0011101; // Expected: {'Z': -1102}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011010; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2564,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011001; Y = 7'b0001001; // Expected: {'Z': -351}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011001; Y = 7'b0001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2565,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -351
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011101; Y = 7'b0010110; // Expected: {'Z': -770}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011101; Y = 7'b0010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2566,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -770
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011010; Y = 7'b1001110; // Expected: {'Z': 1900}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011010; Y = 7'b1001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2567,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101010; Y = 7'b0110010; // Expected: {'Z': 2100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101010; Y = 7'b0110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2568,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b1001011; // Expected: {'Z': -1060}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b1001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2569,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110101; Y = 7'b0110110; // Expected: {'Z': -594}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110101; Y = 7'b0110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2570,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -594
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b0100110; // Expected: {'Z': 342}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2571,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 342
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000111; Y = 7'b0000111; // Expected: {'Z': -399}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000111; Y = 7'b0000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2572,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -399
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001011; Y = 7'b1110110; // Expected: {'Z': 530}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001011; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2573,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 530
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011011; Y = 7'b1010111; // Expected: {'Z': 1517}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011011; Y = 7'b1010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2574,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1517
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b0101101; // Expected: {'Z': -135}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b0101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2575,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110111; Y = 7'b0110111; // Expected: {'Z': 3025}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110111; Y = 7'b0110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2576,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3025
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011001; Y = 7'b0011101; // Expected: {'Z': -1131}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011001; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2577,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b0010010; // Expected: {'Z': 378}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b0010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2578,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 378
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b0001010; // Expected: {'Z': -120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b0001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2579,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110111; Y = 7'b0001000; // Expected: {'Z': -72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110111; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2580,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b0111111; // Expected: {'Z': 3276}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b0111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2581,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3276
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011011; Y = 7'b0100011; // Expected: {'Z': -1295}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011011; Y = 7'b0100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2582,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1295
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011111; Y = 7'b1001000; // Expected: {'Z': -1736}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011111; Y = 7'b1001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2583,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b0000101; // Expected: {'Z': -50}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b0000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2584,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001101; Y = 7'b1000100; // Expected: {'Z': -780}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001101; Y = 7'b1000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2585,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b0110101; // Expected: {'Z': -2226}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2586,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2226
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100010; Y = 7'b1111100; // Expected: {'Z': -136}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100010; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2587,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b1111010; // Expected: {'Z': 168}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b1111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2588,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b1011110; // Expected: {'Z': 612}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b1011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2589,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100001; Y = 7'b0111010; // Expected: {'Z': -1798}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100001; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2590,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101011; Y = 7'b0000010; // Expected: {'Z': -42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101011; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2591,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011010; Y = 7'b1010101; // Expected: {'Z': -1118}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011010; Y = 7'b1010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2592,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001000; Y = 7'b1111101; // Expected: {'Z': -24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001000; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2593,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100111; Y = 7'b1010001; // Expected: {'Z': -1833}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100111; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2594,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1833
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b1101111; // Expected: {'Z': -340}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b1101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2595,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111100; Y = 7'b0011101; // Expected: {'Z': 1740}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111100; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2596,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1740
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101001; Y = 7'b0111111; // Expected: {'Z': 2583}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101001; Y = 7'b0111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2597,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2583
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b0000100; // Expected: {'Z': -192}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b0000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2598,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b0000111; // Expected: {'Z': 119}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b0000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2599,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 119
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101110; Y = 7'b1101001; // Expected: {'Z': -1058}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101110; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2600,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1058
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101011; Y = 7'b1111110; // Expected: {'Z': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101011; Y = 7'b1111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2601,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110101; Y = 7'b1010001; // Expected: {'Z': 517}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110101; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2602,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 517
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100110; Y = 7'b1101100; // Expected: {'Z': 520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100110; Y = 7'b1101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2603,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110001; Y = 7'b1100110; // Expected: {'Z': -1274}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110001; Y = 7'b1100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2604,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1274
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100011; Y = 7'b1101011; // Expected: {'Z': 609}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100011; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2605,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 609
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011101; Y = 7'b1100111; // Expected: {'Z': 875}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011101; Y = 7'b1100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2606,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 875
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b0111101; // Expected: {'Z': -1952}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b0111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2607,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1952
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b1101001; // Expected: {'Z': 1449}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2608,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1449
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111010; Y = 7'b0101011; // Expected: {'Z': 2494}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111010; Y = 7'b0101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2609,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2494
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111100; Y = 7'b0110111; // Expected: {'Z': -220}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111100; Y = 7'b0110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2610,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110111; Y = 7'b0111000; // Expected: {'Z': 3080}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110111; Y = 7'b0111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2611,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100110; Y = 7'b1000101; // Expected: {'Z': 1534}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100110; Y = 7'b1000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2612,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1534
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b1010101; // Expected: {'Z': -731}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b1010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2613,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -731
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b1111010; // Expected: {'Z': -6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b1111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2614,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b0111001; // Expected: {'Z': 2964}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b0111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2615,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2964
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111001; Y = 7'b0100011; // Expected: {'Z': -245}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111001; Y = 7'b0100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2616,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111011; Y = 7'b1000101; // Expected: {'Z': 295}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111011; Y = 7'b1000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2617,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 295
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b1101010; // Expected: {'Z': 880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b1101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2618,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b1001101; // Expected: {'Z': 2448}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b1001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2619,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2448
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b0101001; // Expected: {'Z': -615}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2620,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -615
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111100; Y = 7'b0111011; // Expected: {'Z': 3540}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111100; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2621,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b1000010; // Expected: {'Z': -2790}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b1000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2622,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2790
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100101; Y = 7'b1111100; // Expected: {'Z': -148}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100101; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2623,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b0110100; // Expected: {'Z': -2184}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b0110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2624,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000110; Y = 7'b0010100; // Expected: {'Z': 120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000110; Y = 7'b0010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2625,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011001; Y = 7'b0001110; // Expected: {'Z': -546}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011001; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2626,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b1011010; // Expected: {'Z': 1292}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b1011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2627,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1292
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b1110001; // Expected: {'Z': -45}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b1110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2628,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b1001111; // Expected: {'Z': 1666}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b1001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2629,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1666
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111100; Y = 7'b0001000; // Expected: {'Z': -32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111100; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2630,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111100; Y = 7'b0100100; // Expected: {'Z': -144}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111100; Y = 7'b0100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2631,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001011; Y = 7'b0010110; // Expected: {'Z': -1166}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001011; Y = 7'b0010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2632,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110001; Y = 7'b0101010; // Expected: {'Z': 2058}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110001; Y = 7'b0101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2633,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2058
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000101; Y = 7'b1110001; // Expected: {'Z': -75}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000101; Y = 7'b1110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2634,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011010; Y = 7'b0100110; // Expected: {'Z': -1444}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011010; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2635,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1444
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000000; Y = 7'b1000010; // Expected: {'Z': 3968}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000000; Y = 7'b1000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2636,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3968
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b1010101; // Expected: {'Z': -43}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b1010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2637,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011101; Y = 7'b1111010; // Expected: {'Z': -174}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011101; Y = 7'b1111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2638,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011010; Y = 7'b1101011; // Expected: {'Z': 798}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011010; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2639,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b1110101; // Expected: {'Z': -231}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b1110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2640,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b1101011; // Expected: {'Z': 315}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2641,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 315
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101010; Y = 7'b1100000; // Expected: {'Z': 704}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101010; Y = 7'b1100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2642,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 704
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001010; Y = 7'b0101001; // Expected: {'Z': -2214}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001010; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2643,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101111; Y = 7'b1100110; // Expected: {'Z': -1222}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101111; Y = 7'b1100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2644,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b0111111; // Expected: {'Z': -3024}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b0111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2645,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111100; Y = 7'b1110100; // Expected: {'Z': 48}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111100; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2646,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100100; Y = 7'b0010101; // Expected: {'Z': 756}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100100; Y = 7'b0010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2647,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010110; Y = 7'b1000111; // Expected: {'Z': -1254}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010110; Y = 7'b1000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2648,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000110; Y = 7'b1110000; // Expected: {'Z': 928}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000110; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2649,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 928
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010110; Y = 7'b0101110; // Expected: {'Z': 1012}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010110; Y = 7'b0101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2650,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1012
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b1011110; // Expected: {'Z': 1020}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b1011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2651,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1020
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b1100000; // Expected: {'Z': -1664}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b1100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2652,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1664
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100111; Y = 7'b0010010; // Expected: {'Z': -450}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100111; Y = 7'b0010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2653,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111110; Y = 7'b0100000; // Expected: {'Z': -64}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111110; Y = 7'b0100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2654,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b1011101; // Expected: {'Z': -2170}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b1011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2655,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001100; Y = 7'b0111100; // Expected: {'Z': 720}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001100; Y = 7'b0111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2656,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101000; Y = 7'b0110100; // Expected: {'Z': -1248}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101000; Y = 7'b0110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2657,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100111; Y = 7'b0111100; // Expected: {'Z': -1500}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100111; Y = 7'b0111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2658,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100101; Y = 7'b1001100; // Expected: {'Z': 1404}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100101; Y = 7'b1001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2659,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1404
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001010; Y = 7'b1010101; // Expected: {'Z': -430}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001010; Y = 7'b1010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2660,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b0000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b0000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2661,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b0110111; // Expected: {'Z': -1760}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b0110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2662,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000101; Y = 7'b0100101; // Expected: {'Z': -2183}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000101; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2663,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101001; Y = 7'b0010011; // Expected: {'Z': 779}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101001; Y = 7'b0010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2664,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 779
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000111; Y = 7'b0010001; // Expected: {'Z': -969}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000111; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2665,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -969
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000100; Y = 7'b0011110; // Expected: {'Z': -1800}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000100; Y = 7'b0011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2666,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111111; Y = 7'b1011100; // Expected: {'Z': -2268}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111111; Y = 7'b1011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2667,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2268
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b0000110; // Expected: {'Z': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b0000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2668,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011001; Y = 7'b0010111; // Expected: {'Z': 575}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011001; Y = 7'b0010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2669,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 575
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010110; Y = 7'b0001010; // Expected: {'Z': 220}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010110; Y = 7'b0001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2670,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100111; Y = 7'b1000111; // Expected: {'Z': 1425}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100111; Y = 7'b1000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2671,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1425
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011011; Y = 7'b0100101; // Expected: {'Z': 999}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011011; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2672,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 999
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001000; Y = 7'b0111000; // Expected: {'Z': 448}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001000; Y = 7'b0111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2673,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 448
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000100; Y = 7'b1111101; // Expected: {'Z': 180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000100; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2674,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001001; Y = 7'b0010000; // Expected: {'Z': -880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001001; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2675,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111101; Y = 7'b0001110; // Expected: {'Z': 854}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111101; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2676,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 854
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b0100101; // Expected: {'Z': 888}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2677,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010010; Y = 7'b0100101; // Expected: {'Z': -1702}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010010; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2678,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1702
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000101; Y = 7'b1100000; // Expected: {'Z': -160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000101; Y = 7'b1100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2679,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b0110001; // Expected: {'Z': -1666}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b0110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2680,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1666
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000000; Y = 7'b0010111; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000000; Y = 7'b0010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2681,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100101; Y = 7'b1111110; // Expected: {'Z': 54}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100101; Y = 7'b1111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2682,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100000; Y = 7'b0111000; // Expected: {'Z': 1792}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100000; Y = 7'b0111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2683,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b1001101; // Expected: {'Z': 1173}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b1001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2684,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1173
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000101; Y = 7'b0101110; // Expected: {'Z': -2714}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000101; Y = 7'b0101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2685,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2714
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000111; Y = 7'b1010100; // Expected: {'Z': 2508}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000111; Y = 7'b1010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2686,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2508
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111011; Y = 7'b0010010; // Expected: {'Z': -90}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111011; Y = 7'b0010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2687,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101010; Y = 7'b1100111; // Expected: {'Z': 550}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101010; Y = 7'b1100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2688,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101111; Y = 7'b1001001; // Expected: {'Z': -2585}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101111; Y = 7'b1001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2689,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2585
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b1000110; // Expected: {'Z': -1218}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b1000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2690,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011010; Y = 7'b1010101; // Expected: {'Z': 1634}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011010; Y = 7'b1010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2691,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1634
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b0000100; // Expected: {'Z': -76}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b0000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2692,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100110; Y = 7'b0100011; // Expected: {'Z': 1330}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100110; Y = 7'b0100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2693,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1330
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b0011001; // Expected: {'Z': -450}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b0011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2694,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b0100000; // Expected: {'Z': -320}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b0100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2695,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100110; Y = 7'b0011000; // Expected: {'Z': -624}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100110; Y = 7'b0011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2696,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b0000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b0000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2697,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100111; Y = 7'b0111111; // Expected: {'Z': 2457}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100111; Y = 7'b0111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2698,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2457
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010011; Y = 7'b1110001; // Expected: {'Z': 675}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010011; Y = 7'b1110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2699,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 675
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101011; Y = 7'b1110110; // Expected: {'Z': -430}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101011; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2700,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101100; Y = 7'b1110100; // Expected: {'Z': -528}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101100; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2701,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000101; Y = 7'b1000101; // Expected: {'Z': -295}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000101; Y = 7'b1000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2702,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -295
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001101; Y = 7'b0000011; // Expected: {'Z': -153}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001101; Y = 7'b0000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2703,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -153
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010110; Y = 7'b0000011; // Expected: {'Z': 66}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010110; Y = 7'b0000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2704,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b1110001; // Expected: {'Z': 285}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b1110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2705,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 285
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101111; Y = 7'b0010001; // Expected: {'Z': 799}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101111; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2706,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 799
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100011; Y = 7'b0001100; // Expected: {'Z': -348}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100011; Y = 7'b0001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2707,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -348
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b0100111; // Expected: {'Z': -468}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b0100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2708,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -468
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111000; Y = 7'b1100101; // Expected: {'Z': 216}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111000; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2709,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000110; Y = 7'b1110110; // Expected: {'Z': -60}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000110; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2710,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100000; Y = 7'b0010110; // Expected: {'Z': 704}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100000; Y = 7'b0010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2711,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 704
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001100; Y = 7'b0100101; // Expected: {'Z': -1924}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001100; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2712,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1924
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b1110011; // Expected: {'Z': -117}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2713,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b0011011; // Expected: {'Z': -864}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b0011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2714,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -864
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000101; Y = 7'b1100000; // Expected: {'Z': -160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000101; Y = 7'b1100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2715,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011011; Y = 7'b0011110; // Expected: {'Z': -1110}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011011; Y = 7'b0011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2716,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100101; Y = 7'b1000100; // Expected: {'Z': -2220}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100101; Y = 7'b1000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2717,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b0110010; // Expected: {'Z': -500}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b0110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2718,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b0001000; // Expected: {'Z': -24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2719,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101000; Y = 7'b1001110; // Expected: {'Z': 1200}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101000; Y = 7'b1001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2720,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110110; Y = 7'b1110010; // Expected: {'Z': -756}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110110; Y = 7'b1110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2721,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010000; Y = 7'b0100110; // Expected: {'Z': 608}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010000; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2722,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 608
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010010; Y = 7'b0100101; // Expected: {'Z': 666}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010010; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2723,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 666
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b1110011; // Expected: {'Z': 520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2724,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100111; Y = 7'b1101001; // Expected: {'Z': 575}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100111; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2725,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 575
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b1111001; // Expected: {'Z': 441}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b1111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2726,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 441
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110111; Y = 7'b0111111; // Expected: {'Z': 3465}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110111; Y = 7'b0111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2727,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3465
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011111; Y = 7'b1101001; // Expected: {'Z': -713}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011111; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2728,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -713
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011101; Y = 7'b0100111; // Expected: {'Z': -1365}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011101; Y = 7'b0100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2729,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1365
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b1100010; // Expected: {'Z': 840}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2730,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001101; Y = 7'b0000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001101; Y = 7'b0000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2731,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b1011111; // Expected: {'Z': -2046}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2732,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2046
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110010; Y = 7'b1001111; // Expected: {'Z': 686}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110010; Y = 7'b1001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2733,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 686
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b1000000; // Expected: {'Z': -1344}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b1000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2734,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1344
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000010; Y = 7'b0101111; // Expected: {'Z': 94}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000010; Y = 7'b0101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2735,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010011; Y = 7'b0011011; // Expected: {'Z': 513}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010011; Y = 7'b0011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2736,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 513
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000100; Y = 7'b1100100; // Expected: {'Z': -112}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000100; Y = 7'b1100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2737,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101001; Y = 7'b0000100; // Expected: {'Z': 164}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101001; Y = 7'b0000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2738,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111010; Y = 7'b0001110; // Expected: {'Z': 812}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111010; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2739,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 812
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000100; Y = 7'b1011011; // Expected: {'Z': -148}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000100; Y = 7'b1011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2740,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011100; Y = 7'b1011100; // Expected: {'Z': -1008}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011100; Y = 7'b1011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2741,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b1101011; // Expected: {'Z': 63}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2742,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000101; Y = 7'b1011111; // Expected: {'Z': -165}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000101; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2743,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001000; Y = 7'b1101101; // Expected: {'Z': -152}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001000; Y = 7'b1101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2744,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011101; Y = 7'b1011111; // Expected: {'Z': -957}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011101; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2745,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -957
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101100; Y = 7'b0011101; // Expected: {'Z': 1276}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101100; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2746,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1276
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001100; Y = 7'b1111001; // Expected: {'Z': 364}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001100; Y = 7'b1111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2747,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011100; Y = 7'b1001110; // Expected: {'Z': -1400}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011100; Y = 7'b1001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2748,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000100; Y = 7'b0001111; // Expected: {'Z': 60}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000100; Y = 7'b0001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2749,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001000; Y = 7'b0001101; // Expected: {'Z': 104}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001000; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2750,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b1100110; // Expected: {'Z': -546}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b1100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2751,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101100; Y = 7'b0101001; // Expected: {'Z': 1804}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101100; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2752,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1804
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b0111101; // Expected: {'Z': -2440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b0111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2753,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b0011101; // Expected: {'Z': -1392}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2754,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b0001111; // Expected: {'Z': -450}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b0001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2755,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100011; Y = 7'b1100101; // Expected: {'Z': 783}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100011; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2756,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 783
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001011; Y = 7'b0001110; // Expected: {'Z': -742}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001011; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2757,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -742
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b1000101; // Expected: {'Z': 1770}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b1000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2758,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1770
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010001; Y = 7'b0010101; // Expected: {'Z': -987}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010001; Y = 7'b0010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2759,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -987
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b0001111; // Expected: {'Z': 780}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b0001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2760,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101110; Y = 7'b1011001; // Expected: {'Z': -1794}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101110; Y = 7'b1011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2761,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1794
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100100; Y = 7'b0111111; // Expected: {'Z': 2268}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100100; Y = 7'b0111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2762,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2268
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101010; Y = 7'b1111000; // Expected: {'Z': -336}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101010; Y = 7'b1111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2763,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -336
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111010; Y = 7'b0011100; // Expected: {'Z': -168}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111010; Y = 7'b0011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2764,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100111; Y = 7'b0010000; // Expected: {'Z': 624}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100111; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2765,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b1111101; // Expected: {'Z': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2766,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100111; Y = 7'b1101101; // Expected: {'Z': -741}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100111; Y = 7'b1101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2767,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -741
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101100; Y = 7'b0010001; // Expected: {'Z': 748}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101100; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2768,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 748
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000110; Y = 7'b1011110; // Expected: {'Z': 1972}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000110; Y = 7'b1011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2769,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1972
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b0001000; // Expected: {'Z': -224}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2770,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b0011110; // Expected: {'Z': -570}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b0011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2771,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -570
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100011; Y = 7'b0010011; // Expected: {'Z': -551}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100011; Y = 7'b0010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2772,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -551
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b0101011; // Expected: {'Z': -731}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b0101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2773,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -731
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111010; Y = 7'b0110110; // Expected: {'Z': 3132}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111010; Y = 7'b0110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2774,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b1101101; // Expected: {'Z': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b1101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2775,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111100; Y = 7'b1000000; // Expected: {'Z': 256}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111100; Y = 7'b1000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2776,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 256
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010011; Y = 7'b0011101; // Expected: {'Z': -1305}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010011; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2777,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1305
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001100; Y = 7'b0001110; // Expected: {'Z': 168}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001100; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2778,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001110; Y = 7'b0110101; // Expected: {'Z': 742}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001110; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2779,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 742
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001100; Y = 7'b1001101; // Expected: {'Z': -612}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001100; Y = 7'b1001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2780,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000101; Y = 7'b1111001; // Expected: {'Z': -35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000101; Y = 7'b1111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2781,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b1100010; // Expected: {'Z': -1560}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b1100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2782,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111101; Y = 7'b1110110; // Expected: {'Z': -610}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111101; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2783,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -610
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b1100011; // Expected: {'Z': 435}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b1100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2784,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 435
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110011; Y = 7'b1010111; // Expected: {'Z': -2091}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110011; Y = 7'b1010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2785,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2091
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b0010011; // Expected: {'Z': -912}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b0010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2786,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -912
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b0000111; // Expected: {'Z': -7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b0000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2787,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b1101111; // Expected: {'Z': 680}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b1101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2788,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100010; Y = 7'b0001001; // Expected: {'Z': 306}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100010; Y = 7'b0001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2789,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 306
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001100; Y = 7'b0101011; // Expected: {'Z': -2236}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001100; Y = 7'b0101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2790,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110000; Y = 7'b0110001; // Expected: {'Z': -784}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110000; Y = 7'b0110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2791,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100111; Y = 7'b0110110; // Expected: {'Z': 2106}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100111; Y = 7'b0110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2792,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000110; Y = 7'b0000110; // Expected: {'Z': 36}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000110; Y = 7'b0000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2793,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100001; Y = 7'b0111011; // Expected: {'Z': 1947}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100001; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2794,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1947
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101110; Y = 7'b1100011; // Expected: {'Z': -1334}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101110; Y = 7'b1100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2795,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1334
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b0000001; // Expected: {'Z': -42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b0000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2796,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b0001000; // Expected: {'Z': -240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2797,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b0000110; // Expected: {'Z': 54}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b0000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2798,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001010; Y = 7'b1000000; // Expected: {'Z': 3456}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001010; Y = 7'b1000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2799,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010000; Y = 7'b1110100; // Expected: {'Z': 576}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010000; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2800,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b0101110; // Expected: {'Z': 920}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b0101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2801,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110000; Y = 7'b1111001; // Expected: {'Z': 112}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110000; Y = 7'b1111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2802,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011100; Y = 7'b0111000; // Expected: {'Z': 1568}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011100; Y = 7'b0111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2803,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1568
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110010; Y = 7'b1110011; // Expected: {'Z': -650}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110010; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2804,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011001; Y = 7'b1010111; // Expected: {'Z': 1599}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011001; Y = 7'b1010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2805,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1599
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011100; Y = 7'b0000001; // Expected: {'Z': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011100; Y = 7'b0000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2806,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010000; Y = 7'b1110110; // Expected: {'Z': -160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010000; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2807,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001010; Y = 7'b1101100; // Expected: {'Z': 1080}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001010; Y = 7'b1101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2808,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011111; Y = 7'b1101101; // Expected: {'Z': 627}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011111; Y = 7'b1101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2809,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 627
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b1011000; // Expected: {'Z': 920}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b1011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2810,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111000; Y = 7'b1111011; // Expected: {'Z': -280}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111000; Y = 7'b1111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2811,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100110; Y = 7'b1110001; // Expected: {'Z': -570}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100110; Y = 7'b1110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2812,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -570
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001111; Y = 7'b1001111; // Expected: {'Z': -735}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001111; Y = 7'b1001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2813,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -735
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001101; Y = 7'b1111100; // Expected: {'Z': -52}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001101; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2814,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111110; Y = 7'b1000000; // Expected: {'Z': 128}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111110; Y = 7'b1000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2815,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011101; Y = 7'b0000111; // Expected: {'Z': 203}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011101; Y = 7'b0000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2816,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 203
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000000; Y = 7'b1001100; // Expected: {'Z': 3328}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000000; Y = 7'b1001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2817,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3328
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111001; Y = 7'b0110001; // Expected: {'Z': 2793}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111001; Y = 7'b0110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2818,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2793
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100101; Y = 7'b1011111; // Expected: {'Z': 891}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100101; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2819,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 891
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010001; Y = 7'b0001000; // Expected: {'Z': -376}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010001; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2820,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -376
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b1010001; // Expected: {'Z': -423}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2821,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -423
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111101; Y = 7'b1101111; // Expected: {'Z': -1037}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111101; Y = 7'b1101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2822,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1037
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001111; Y = 7'b0000100; // Expected: {'Z': -196}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001111; Y = 7'b0000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2823,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101000; Y = 7'b1010100; // Expected: {'Z': 1056}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101000; Y = 7'b1010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2824,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1056
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101011; Y = 7'b0100111; // Expected: {'Z': -819}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101011; Y = 7'b0100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2825,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -819
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b1110101; // Expected: {'Z': -572}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b1110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2826,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -572
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111010; Y = 7'b1011010; // Expected: {'Z': -2204}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111010; Y = 7'b1011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2827,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100001; Y = 7'b1111100; // Expected: {'Z': 124}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100001; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2828,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b1101000; // Expected: {'Z': 480}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b1101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2829,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b0010010; // Expected: {'Z': -414}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b0010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2830,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -414
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111000; Y = 7'b0011101; // Expected: {'Z': -232}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111000; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2831,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000111; Y = 7'b0110111; // Expected: {'Z': 385}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000111; Y = 7'b0110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2832,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 385
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100111; Y = 7'b1111111; // Expected: {'Z': -39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100111; Y = 7'b1111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2833,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111001; Y = 7'b0110101; // Expected: {'Z': 3021}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111001; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2834,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3021
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b1101011; // Expected: {'Z': 483}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2835,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 483
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010111; Y = 7'b1011001; // Expected: {'Z': 1599}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010111; Y = 7'b1011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2836,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1599
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011101; Y = 7'b0011011; // Expected: {'Z': 783}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011101; Y = 7'b0011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2837,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 783
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b1111110; // Expected: {'Z': 126}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b1111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2838,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110000; Y = 7'b0001100; // Expected: {'Z': -192}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110000; Y = 7'b0001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2839,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110011; Y = 7'b1001011; // Expected: {'Z': -2703}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110011; Y = 7'b1001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2840,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2703
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b0110011; // Expected: {'Z': -3213}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b0110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2841,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b0010110; // Expected: {'Z': -330}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b0010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2842,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -330
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111010; Y = 7'b1110100; // Expected: {'Z': 72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111010; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2843,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b1011011; // Expected: {'Z': 740}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b1011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2844,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 740
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001001; Y = 7'b0111010; // Expected: {'Z': -3190}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001001; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2845,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001000; Y = 7'b1001110; // Expected: {'Z': 2800}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001000; Y = 7'b1001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2846,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b1001011; // Expected: {'Z': 1590}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b1001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2847,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1590
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111100; Y = 7'b0001101; // Expected: {'Z': -52}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111100; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2848,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011010; Y = 7'b0110011; // Expected: {'Z': -1938}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011010; Y = 7'b0110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2849,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1938
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100011; Y = 7'b0110101; // Expected: {'Z': 1855}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100011; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2850,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1855
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110111; Y = 7'b0110100; // Expected: {'Z': -468}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110111; Y = 7'b0110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2851,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -468
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110000; Y = 7'b0011110; // Expected: {'Z': -480}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110000; Y = 7'b0011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2852,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100101; Y = 7'b1010000; // Expected: {'Z': 1296}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100101; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2853,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010011; Y = 7'b0100111; // Expected: {'Z': -1755}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010011; Y = 7'b0100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2854,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1755
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b1001101; // Expected: {'Z': -51}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b1001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2855,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111101; Y = 7'b0000011; // Expected: {'Z': 183}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111101; Y = 7'b0000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2856,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100101; Y = 7'b1010100; // Expected: {'Z': 1188}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100101; Y = 7'b1010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2857,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b0001100; // Expected: {'Z': 744}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b0001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2858,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 744
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111001; Y = 7'b1010011; // Expected: {'Z': 315}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111001; Y = 7'b1010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2859,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 315
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b1010000; // Expected: {'Z': 1440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2860,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110010; Y = 7'b0001110; // Expected: {'Z': -196}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110010; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2861,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b1011110; // Expected: {'Z': 1428}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b1011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2862,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1428
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b0001001; // Expected: {'Z': -135}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b0001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2863,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110110; Y = 7'b1100011; // Expected: {'Z': -1566}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110110; Y = 7'b1100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2864,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1566
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010010; Y = 7'b0010000; // Expected: {'Z': 288}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010010; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2865,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110101; Y = 7'b0110101; // Expected: {'Z': -583}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110101; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2866,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -583
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110001; Y = 7'b1110000; // Expected: {'Z': -784}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110001; Y = 7'b1110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2867,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011110; Y = 7'b1101011; // Expected: {'Z': -630}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011110; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2868,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -630
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011011; Y = 7'b1011100; // Expected: {'Z': 1332}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011011; Y = 7'b1011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2869,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1332
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000100; Y = 7'b0111111; // Expected: {'Z': 252}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000100; Y = 7'b0111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2870,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b1110101; // Expected: {'Z': -33}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b1110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2871,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001111; Y = 7'b1111000; // Expected: {'Z': 392}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001111; Y = 7'b1111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2872,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111001; Y = 7'b0011111; // Expected: {'Z': -217}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111001; Y = 7'b0011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2873,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111011; Y = 7'b0110010; // Expected: {'Z': 2950}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111011; Y = 7'b0110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2874,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011010; Y = 7'b0100110; // Expected: {'Z': -1444}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011010; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2875,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1444
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111000; Y = 7'b0011111; // Expected: {'Z': -248}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111000; Y = 7'b0011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2876,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100011; Y = 7'b1001100; // Expected: {'Z': -1820}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100011; Y = 7'b1001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2877,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b1101000; // Expected: {'Z': -24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b1101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2878,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b1101000; // Expected: {'Z': 360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b1101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2879,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111110; Y = 7'b0000101; // Expected: {'Z': -10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111110; Y = 7'b0000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2880,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000101; Y = 7'b1011101; // Expected: {'Z': 2065}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000101; Y = 7'b1011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2881,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2065
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001110; Y = 7'b0100111; // Expected: {'Z': 546}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001110; Y = 7'b0100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2882,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b1111101; // Expected: {'Z': 108}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2883,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b0101011; // Expected: {'Z': 2279}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b0101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2884,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2279
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101010; Y = 7'b1110110; // Expected: {'Z': -420}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101010; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2885,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101000; Y = 7'b1000001; // Expected: {'Z': 1512}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101000; Y = 7'b1000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2886,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1512
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b0001001; // Expected: {'Z': -9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b0001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2887,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101001; Y = 7'b0000111; // Expected: {'Z': 287}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101001; Y = 7'b0000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2888,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 287
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010110; Y = 7'b1000101; // Expected: {'Z': 2478}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010110; Y = 7'b1000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2889,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2478
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b1001111; // Expected: {'Z': 490}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b1001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2890,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 490
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110011; Y = 7'b1010110; // Expected: {'Z': 546}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110011; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2891,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000000; Y = 7'b1101001; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000000; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2892,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b0011000; // Expected: {'Z': -480}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b0011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2893,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111100; Y = 7'b1100111; // Expected: {'Z': -1500}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111100; Y = 7'b1100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2894,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100111; Y = 7'b0101101; // Expected: {'Z': -1125}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100111; Y = 7'b0101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2895,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011111; Y = 7'b1000100; // Expected: {'Z': 1980}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011111; Y = 7'b1000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2896,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b0101100; // Expected: {'Z': -1232}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b0101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2897,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011111; Y = 7'b1010110; // Expected: {'Z': 1386}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011111; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2898,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1386
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100001; Y = 7'b1001000; // Expected: {'Z': -1848}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100001; Y = 7'b1001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2899,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010010; Y = 7'b0111011; // Expected: {'Z': -2714}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010010; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2900,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2714
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b0010000; // Expected: {'Z': 320}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2901,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b0010110; // Expected: {'Z': -66}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b0010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2902,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001000; Y = 7'b1000111; // Expected: {'Z': -456}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001000; Y = 7'b1000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2903,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011001; Y = 7'b1011110; // Expected: {'Z': 1326}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011001; Y = 7'b1011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2904,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1326
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000101; Y = 7'b1111100; // Expected: {'Z': -20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000101; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2905,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010101; Y = 7'b1001000; // Expected: {'Z': 2408}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010101; Y = 7'b1001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2906,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011010; Y = 7'b1000110; // Expected: {'Z': -1508}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011010; Y = 7'b1000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2907,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1508
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111001; Y = 7'b0001110; // Expected: {'Z': 798}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111001; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2908,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b1001100; // Expected: {'Z': 1456}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b1001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2909,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100011; Y = 7'b1000000; // Expected: {'Z': -2240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100011; Y = 7'b1000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2910,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010100; Y = 7'b1011100; // Expected: {'Z': -720}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010100; Y = 7'b1011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2911,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001101; Y = 7'b0110001; // Expected: {'Z': 637}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001101; Y = 7'b0110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2912,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 637
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000110; Y = 7'b1000100; // Expected: {'Z': 3480}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000110; Y = 7'b1000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2913,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111110; Y = 7'b0011111; // Expected: {'Z': 1922}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111110; Y = 7'b0011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2914,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1922
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111010; Y = 7'b1100000; // Expected: {'Z': -1856}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111010; Y = 7'b1100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2915,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000011; Y = 7'b1001110; // Expected: {'Z': 3050}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000011; Y = 7'b1001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2916,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110101; Y = 7'b1001010; // Expected: {'Z': 594}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110101; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2917,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 594
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000010; Y = 7'b1110111; // Expected: {'Z': -18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000010; Y = 7'b1110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2918,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b1100100; // Expected: {'Z': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b1100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2919,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110011; Y = 7'b1111111; // Expected: {'Z': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110011; Y = 7'b1111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2920,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001110; Y = 7'b0001110; // Expected: {'Z': 196}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001110; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2921,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010010; Y = 7'b1001011; // Expected: {'Z': -954}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010010; Y = 7'b1001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2922,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -954
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001100; Y = 7'b1100011; // Expected: {'Z': -348}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001100; Y = 7'b1100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2923,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -348
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b1111100; // Expected: {'Z': -36}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2924,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b1001111; // Expected: {'Z': 980}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b1001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2925,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b1111101; // Expected: {'Z': 189}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2926,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111110; Y = 7'b0010101; // Expected: {'Z': -42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111110; Y = 7'b0010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2927,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101001; Y = 7'b1001101; // Expected: {'Z': -2091}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101001; Y = 7'b1001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2928,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2091
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b0000011; // Expected: {'Z': -108}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b0000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2929,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b0010111; // Expected: {'Z': -391}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b0010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2930,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -391
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000010; Y = 7'b1101000; // Expected: {'Z': 1488}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000010; Y = 7'b1101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2931,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101010; Y = 7'b1000101; // Expected: {'Z': 1298}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101010; Y = 7'b1000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2932,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1298
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101101; Y = 7'b1101011; // Expected: {'Z': 399}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101101; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2933,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 399
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100000; Y = 7'b0010111; // Expected: {'Z': -736}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100000; Y = 7'b0010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2934,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011110; Y = 7'b0101001; // Expected: {'Z': -1394}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011110; Y = 7'b0101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2935,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1394
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b1010100; // Expected: {'Z': -1056}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b1010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2936,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1056
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111101; Y = 7'b1111000; // Expected: {'Z': -488}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111101; Y = 7'b1111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2937,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b1100110; // Expected: {'Z': -442}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b1100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2938,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -442
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100110; Y = 7'b1010110; // Expected: {'Z': -1596}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100110; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2939,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1596
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111010; Y = 7'b0101110; // Expected: {'Z': 2668}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111010; Y = 7'b0101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2940,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2668
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000111; Y = 7'b1011111; // Expected: {'Z': -231}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000111; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2941,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000101; Y = 7'b0010001; // Expected: {'Z': 85}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000101; Y = 7'b0010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2942,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 85
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011011; Y = 7'b1010100; // Expected: {'Z': 1628}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011011; Y = 7'b1010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2943,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1628
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b1000000; // Expected: {'Z': -2880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b1000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2944,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100001; Y = 7'b0000011; // Expected: {'Z': 99}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100001; Y = 7'b0000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2945,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000011; Y = 7'b1001010; // Expected: {'Z': 3294}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000011; Y = 7'b1001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2946,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3294
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110000; Y = 7'b0100110; // Expected: {'Z': -608}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110000; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2947,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -608
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010111; Y = 7'b0010000; // Expected: {'Z': -656}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010111; Y = 7'b0010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2948,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -656
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b0001101; // Expected: {'Z': -520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2949,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100101; Y = 7'b0000110; // Expected: {'Z': 222}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100101; Y = 7'b0000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2950,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110101; Y = 7'b1100111; // Expected: {'Z': 275}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110101; Y = 7'b1100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2951,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 275
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101001; Y = 7'b0001001; // Expected: {'Z': 369}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101001; Y = 7'b0001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2952,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 369
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b0010101; // Expected: {'Z': -63}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b0010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2953,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000100; Y = 7'b1100100; // Expected: {'Z': 1680}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000100; Y = 7'b1100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2954,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111111; Y = 7'b0001001; // Expected: {'Z': 567}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111111; Y = 7'b0001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2955,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 567
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111011; Y = 7'b1101101; // Expected: {'Z': 95}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111011; Y = 7'b1101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2956,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b1011011; // Expected: {'Z': -111}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b1011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2957,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -111
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000100; Y = 7'b0010110; // Expected: {'Z': -1320}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000100; Y = 7'b0010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2958,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011010; Y = 7'b0011100; // Expected: {'Z': 728}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011010; Y = 7'b0011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2959,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011001; Y = 7'b0011110; // Expected: {'Z': 750}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011001; Y = 7'b0011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2960,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101011; Y = 7'b0100100; // Expected: {'Z': 1548}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101011; Y = 7'b0100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2961,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1548
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010010; Y = 7'b0101111; // Expected: {'Z': 846}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010010; Y = 7'b0101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2962,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 846
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011100; Y = 7'b0100101; // Expected: {'Z': 1036}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011100; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2963,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1036
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101011; Y = 7'b1110001; // Expected: {'Z': -645}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101011; Y = 7'b1110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2964,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -645
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b1000000; // Expected: {'Z': 1792}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b1000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2965,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011111; Y = 7'b0101110; // Expected: {'Z': -1518}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011111; Y = 7'b0101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2966,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1518
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100011; Y = 7'b0100110; // Expected: {'Z': -1102}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100011; Y = 7'b0100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2967,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001010; Y = 7'b0100000; // Expected: {'Z': 320}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001010; Y = 7'b0100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2968,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010100; Y = 7'b0001101; // Expected: {'Z': -572}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010100; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2969,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -572
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b0100010; // Expected: {'Z': -2142}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b0100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2970,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011001; Y = 7'b0000100; // Expected: {'Z': 100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011001; Y = 7'b0000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2971,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011001; Y = 7'b0110010; // Expected: {'Z': 1250}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011001; Y = 7'b0110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2972,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100101; Y = 7'b1011111; // Expected: {'Z': -1221}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100101; Y = 7'b1011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2973,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110111; Y = 7'b0001010; // Expected: {'Z': 550}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110111; Y = 7'b0001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2974,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b1001111; // Expected: {'Z': -147}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b1001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2975,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b1010010; // Expected: {'Z': 690}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b1010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2976,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 690
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001110; Y = 7'b1000100; // Expected: {'Z': -840}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001110; Y = 7'b1000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2977,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001010; Y = 7'b1111100; // Expected: {'Z': 216}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001010; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2978,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111101; Y = 7'b1111001; // Expected: {'Z': -427}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111101; Y = 7'b1111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2979,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -427
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111011; Y = 7'b0001101; // Expected: {'Z': 767}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111011; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2980,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 767
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010000; Y = 7'b1011001; // Expected: {'Z': -624}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010000; Y = 7'b1011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2981,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011000; Y = 7'b0011101; // Expected: {'Z': -1160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011000; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2982,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b1010010; // Expected: {'Z': -2392}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b1010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2983,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101000; Y = 7'b0111011; // Expected: {'Z': -1416}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101000; Y = 7'b0111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2984,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110111; Y = 7'b1001011; // Expected: {'Z': -2915}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110111; Y = 7'b1001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2985,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2915
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b0000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b0000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2986,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001101; Y = 7'b1101100; // Expected: {'Z': -260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001101; Y = 7'b1101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2987,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b0100000; // Expected: {'Z': 544}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b0100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2988,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 544
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b1110110; // Expected: {'Z': -240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2989,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001011; Y = 7'b1111100; // Expected: {'Z': -44}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001011; Y = 7'b1111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2990,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001101; Y = 7'b1100100; // Expected: {'Z': -364}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001101; Y = 7'b1100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2991,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011001; Y = 7'b0110011; // Expected: {'Z': 1275}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011001; Y = 7'b0110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2992,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1275
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100001; Y = 7'b0111100; // Expected: {'Z': 1980}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100001; Y = 7'b0111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2993,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000000; Y = 7'b0010110; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000000; Y = 7'b0010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2994,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101110; Y = 7'b1101111; // Expected: {'Z': -782}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101110; Y = 7'b1101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2995,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -782
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001010; Y = 7'b1101111; // Expected: {'Z': -170}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001010; Y = 7'b1101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2996,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b1100101; // Expected: {'Z': -243}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b1100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2997,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000100; Y = 7'b1111111; // Expected: {'Z': -4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000100; Y = 7'b1111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2998,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011010; Y = 7'b0111001; // Expected: {'Z': 1482}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011010; Y = 7'b0111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2999,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1482
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001010; Y = 7'b0011001; // Expected: {'Z': 250}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001010; Y = 7'b0011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3000,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110000; Y = 7'b1010111; // Expected: {'Z': 656}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110000; Y = 7'b1010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3001,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 656
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b0111111; // Expected: {'Z': 3276}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b0111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3002,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3276
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111100; Y = 7'b1100100; // Expected: {'Z': 112}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111100; Y = 7'b1100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3003,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111100; Y = 7'b1000110; // Expected: {'Z': 232}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111100; Y = 7'b1000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3004,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100000; Y = 7'b0001010; // Expected: {'Z': 320}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100000; Y = 7'b0001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3005,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b0001011; // Expected: {'Z': -187}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b0001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3006,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001100; Y = 7'b0111101; // Expected: {'Z': 732}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001100; Y = 7'b0111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3007,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 732
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111101; Y = 7'b1010000; // Expected: {'Z': -2928}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111101; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3008,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2928
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011110; Y = 7'b1000111; // Expected: {'Z': -1710}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011110; Y = 7'b1000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3009,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1710
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000010; Y = 7'b0011101; // Expected: {'Z': 58}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000010; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3010,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011010; Y = 7'b1101101; // Expected: {'Z': -494}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011010; Y = 7'b1101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3011,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -494
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000010; Y = 7'b1011000; // Expected: {'Z': -80}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000010; Y = 7'b1011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3012,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b0101000; // Expected: {'Z': -1200}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b0101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3013,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110000; Y = 7'b1111010; // Expected: {'Z': -288}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110000; Y = 7'b1111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3014,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000001; Y = 7'b0001011; // Expected: {'Z': -693}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000001; Y = 7'b0001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3015,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -693
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011100; Y = 7'b1101001; // Expected: {'Z': 828}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011100; Y = 7'b1101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3016,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111010; Y = 7'b0011111; // Expected: {'Z': 1798}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111010; Y = 7'b0011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3017,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001111; Y = 7'b0011011; // Expected: {'Z': 405}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001111; Y = 7'b0011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3018,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 405
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b1101011; // Expected: {'Z': 483}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3019,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 483
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001111; Y = 7'b0110101; // Expected: {'Z': -2597}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001111; Y = 7'b0110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3020,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2597
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001011; Y = 7'b0011110; // Expected: {'Z': -1590}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001011; Y = 7'b0011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3021,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1590
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001101; Y = 7'b0001011; // Expected: {'Z': -561}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001101; Y = 7'b0001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3022,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -561
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111011; Y = 7'b0110011; // Expected: {'Z': 3009}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111011; Y = 7'b0110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3023,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3009
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100011; Y = 7'b0111111; // Expected: {'Z': 2205}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100011; Y = 7'b0111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3024,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101000; Y = 7'b0101110; // Expected: {'Z': 1840}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101000; Y = 7'b0101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3025,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100111; Y = 7'b0001100; // Expected: {'Z': -300}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100111; Y = 7'b0001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3026,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000000; Y = 7'b1101011; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000000; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3027,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b1110110; // Expected: {'Z': 230}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3028,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110101; Y = 7'b1010011; // Expected: {'Z': 495}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110101; Y = 7'b1010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3029,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 495
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010011; Y = 7'b1001001; // Expected: {'Z': 2475}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010011; Y = 7'b1001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3030,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2475
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001111; Y = 7'b1010110; // Expected: {'Z': -630}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001111; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3031,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -630
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111010; Y = 7'b1110101; // Expected: {'Z': -638}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111010; Y = 7'b1110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3032,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -638
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111010; Y = 7'b0010100; // Expected: {'Z': -120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111010; Y = 7'b0010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3033,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110011; Y = 7'b1111000; // Expected: {'Z': 104}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110011; Y = 7'b1111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3034,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b1111101; // Expected: {'Z': -9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3035,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011111; Y = 7'b0110010; // Expected: {'Z': 1550}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011111; Y = 7'b0110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3036,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000101; Y = 7'b1000000; // Expected: {'Z': 3776}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000101; Y = 7'b1000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3037,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3776
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101001; Y = 7'b0101100; // Expected: {'Z': 1804}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101001; Y = 7'b0101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3038,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1804
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101101; Y = 7'b0100001; // Expected: {'Z': 1485}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101101; Y = 7'b0100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3039,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1485
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010011; Y = 7'b1111111; // Expected: {'Z': 45}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010011; Y = 7'b1111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3040,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000110; Y = 7'b0000010; // Expected: {'Z': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000110; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3041,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b1111000; // Expected: {'Z': 136}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b1111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3042,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001001; Y = 7'b0001001; // Expected: {'Z': -495}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001001; Y = 7'b0001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3043,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -495
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000011; Y = 7'b1100111; // Expected: {'Z': -75}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000011; Y = 7'b1100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3044,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001100; Y = 7'b0000100; // Expected: {'Z': -208}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001100; Y = 7'b0000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3045,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b1101010; // Expected: {'Z': -462}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b1101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3046,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b0100111; // Expected: {'Z': -780}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b0100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3047,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110011; Y = 7'b0010011; // Expected: {'Z': -247}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110011; Y = 7'b0010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3048,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011011; Y = 7'b1011000; // Expected: {'Z': 1480}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011011; Y = 7'b1011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3049,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110000; Y = 7'b0000101; // Expected: {'Z': -80}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110000; Y = 7'b0000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3050,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111011; Y = 7'b1100100; // Expected: {'Z': -1652}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111011; Y = 7'b1100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3051,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1652
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b1100000; // Expected: {'Z': 384}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b1100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3052,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 384
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000001; Y = 7'b0011000; // Expected: {'Z': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000001; Y = 7'b0011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3053,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b0111110; // Expected: {'Z': -1116}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b0111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3054,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010101; Y = 7'b1110110; // Expected: {'Z': -210}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010101; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3055,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001110; Y = 7'b0010010; // Expected: {'Z': -900}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001110; Y = 7'b0010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3056,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110110; Y = 7'b0100000; // Expected: {'Z': 1728}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110110; Y = 7'b0100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3057,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000110; Y = 7'b1000001; // Expected: {'Z': 3654}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000110; Y = 7'b1000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3058,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3654
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100101; Y = 7'b0111010; // Expected: {'Z': -1566}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100101; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3059,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1566
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101111; Y = 7'b0111101; // Expected: {'Z': -1037}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101111; Y = 7'b0111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3060,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1037
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110011; Y = 7'b1010000; // Expected: {'Z': 624}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110011; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3061,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101001; Y = 7'b1111010; // Expected: {'Z': 138}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101001; Y = 7'b1111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3062,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101000; Y = 7'b1110100; // Expected: {'Z': 288}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101000; Y = 7'b1110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3063,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111001; Y = 7'b0100111; // Expected: {'Z': -273}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111001; Y = 7'b0100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3064,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -273
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100011; Y = 7'b0010100; // Expected: {'Z': -580}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100011; Y = 7'b0010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3065,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b1001100; // Expected: {'Z': 780}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b1001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3066,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101110; Y = 7'b0101000; // Expected: {'Z': -720}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101110; Y = 7'b0101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3067,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011100; Y = 7'b1001011; // Expected: {'Z': -1484}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011100; Y = 7'b1001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3068,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1484
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b1110101; // Expected: {'Z': -583}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b1110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3069,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -583
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101100; Y = 7'b0011000; // Expected: {'Z': 1056}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101100; Y = 7'b0011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3070,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1056
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b1000011; // Expected: {'Z': 61}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b1000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3071,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111100; Y = 7'b0110100; // Expected: {'Z': 3120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111100; Y = 7'b0110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3072,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101000; Y = 7'b1101011; // Expected: {'Z': 504}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101000; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3073,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110101; Y = 7'b0010110; // Expected: {'Z': -242}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110101; Y = 7'b0010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3074,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110011; Y = 7'b1011011; // Expected: {'Z': -1887}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110011; Y = 7'b1011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3075,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1887
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110101; Y = 7'b0000010; // Expected: {'Z': 106}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110101; Y = 7'b0000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3076,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001000; Y = 7'b0001000; // Expected: {'Z': 64}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001000; Y = 7'b0001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3077,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110110; Y = 7'b1110011; // Expected: {'Z': -702}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110110; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3078,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -702
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011010; Y = 7'b1101100; // Expected: {'Z': 760}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011010; Y = 7'b1101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3079,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010111; Y = 7'b1000100; // Expected: {'Z': -1380}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010111; Y = 7'b1000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3080,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1380
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100001; Y = 7'b1010001; // Expected: {'Z': 1457}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100001; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3081,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1457
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100001; Y = 7'b1101011; // Expected: {'Z': 651}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100001; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3082,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 651
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001111; Y = 7'b0111101; // Expected: {'Z': 915}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001111; Y = 7'b0111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3083,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 915
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100010; Y = 7'b0100000; // Expected: {'Z': 1088}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100010; Y = 7'b0100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3084,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1088
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100010; Y = 7'b1111111; // Expected: {'Z': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100010; Y = 7'b1111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3085,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101010; Y = 7'b1011001; // Expected: {'Z': -1638}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101010; Y = 7'b1011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3086,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1638
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b1011101; // Expected: {'Z': -840}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b1011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3087,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100111; Y = 7'b0110011; // Expected: {'Z': -1275}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100111; Y = 7'b0110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3088,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1275
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111011; Y = 7'b1000110; // Expected: {'Z': 290}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111011; Y = 7'b1000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3089,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 290
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011000; Y = 7'b1101011; // Expected: {'Z': -504}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011000; Y = 7'b1101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3090,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0111100; Y = 7'b1001001; // Expected: {'Z': -3300}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0111100; Y = 7'b1001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3091,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101100; Y = 7'b1111010; // Expected: {'Z': 120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101100; Y = 7'b1111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3092,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0000010; Y = 7'b0101011; // Expected: {'Z': 86}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0000010; Y = 7'b0101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3093,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100101; Y = 7'b1110011; // Expected: {'Z': 351}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100101; Y = 7'b1110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3094,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 351
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0001001; Y = 7'b0100101; // Expected: {'Z': 333}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0001001; Y = 7'b0100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3095,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 333
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100110; Y = 7'b0000111; // Expected: {'Z': -182}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100110; Y = 7'b0000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3096,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110110; Y = 7'b0010100; // Expected: {'Z': -200}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110110; Y = 7'b0010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3097,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011011; Y = 7'b0011100; // Expected: {'Z': 756}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011011; Y = 7'b0011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3098,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1011011; Y = 7'b0001110; // Expected: {'Z': -518}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1011011; Y = 7'b0001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3099,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -518
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010011; Y = 7'b0001010; // Expected: {'Z': 190}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010011; Y = 7'b0001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3100,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111111; Y = 7'b1010001; // Expected: {'Z': 47}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111111; Y = 7'b1010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3101,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000000; Y = 7'b0111010; // Expected: {'Z': -3712}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000000; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3102,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3712
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110111; Y = 7'b0001101; // Expected: {'Z': -117}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110111; Y = 7'b0001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3103,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110010; Y = 7'b1010010; // Expected: {'Z': -2300}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110010; Y = 7'b1010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3104,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1010010; Y = 7'b0110100; // Expected: {'Z': -2392}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1010010; Y = 7'b0110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3105,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0010001; Y = 7'b1000101; // Expected: {'Z': -1003}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0010001; Y = 7'b1000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3106,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1003
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100100; Y = 7'b0111010; // Expected: {'Z': -1624}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100100; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3107,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001001; Y = 7'b0011101; // Expected: {'Z': -1595}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001001; Y = 7'b0011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3108,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1595
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0100010; Y = 7'b1010000; // Expected: {'Z': -1632}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0100010; Y = 7'b1010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3109,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1632
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0011011; Y = 7'b1001001; // Expected: {'Z': -1485}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0011011; Y = 7'b1001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3110,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1485
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1111101; Y = 7'b0111111; // Expected: {'Z': -189}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1111101; Y = 7'b0111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3111,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1000100; Y = 7'b0110000; // Expected: {'Z': -2880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1000100; Y = 7'b0110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3112,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1100101; Y = 7'b1010110; // Expected: {'Z': 1134}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1100101; Y = 7'b1010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3113,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b0100000; // Expected: {'Z': 1664}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b0100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3114,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1664
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110001; Y = 7'b1011000; // Expected: {'Z': 600}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110001; Y = 7'b1011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3115,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110111; Y = 7'b0000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110111; Y = 7'b0000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3116,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1101011; Y = 7'b1010011; // Expected: {'Z': 945}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1101011; Y = 7'b1010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3117,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 945
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0110100; Y = 7'b1110110; // Expected: {'Z': -520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0110100; Y = 7'b1110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3118,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1110100; Y = 7'b1111101; // Expected: {'Z': 36}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1110100; Y = 7'b1111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3119,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b1001000; Y = 7'b1011010; // Expected: {'Z': 2128}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b1001000; Y = 7'b1011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3120,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 7'b0101111; Y = 7'b0111010; // Expected: {'Z': 2726}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 7'b0101111; Y = 7'b0111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3121,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2726
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        $finish;
    end
  
endmodule