
`timescale 1ns / 1ps

module tb_N5_restoring_divider;

    // Parameters
    
    parameter N = 5;
    
     
    // Inputs
    
    reg   clk;
    
    reg   rst;
    
    reg   start;
    
    reg  [4:0] X;
    
    reg  [4:0] Y;
    
    
    // Outputs
    
    wire  [4:0] quot;
    
    wire  [4:0] rem;
    
    wire   valid;
    
    
    // Instantiate the Unit Under Test (UUT)
    restoring_divider  #( N ) uut (
        
        .clk(clk),
        
        .rst(rst),
        
        .start(start),
        
        .X(X),
        
        .Y(Y),
        
        
        .quot(quot),
        
        .rem(rem),
        
        .valid(valid)
        
    );

    // Clock generation 
    
    
            always begin
                #5 clk = ~clk;
            end
            
    

    
    
            always begin
                #99 rst = 1'b1; 
            end
            
    
    
    initial begin
        // Initialize Inputs
        
        clk = 0;
        
        rst = 0;
        
        start = 0;
        
        X = 0;
        
        Y = 0;
        
    
        // Wait for global reset
        #100;
    
        // Stimuli
        
        #10 X = 5'b10001; Y = 5'b01111; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 0,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b00011; // Expected: {'quot': 9, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 9, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b11000; // Expected: {'quot': 0, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b11000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 3,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00100; Y = 5'b00100; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00100; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 4,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b01110; // Expected: {'quot': 1, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 5,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b01001; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 6,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11011; Y = 5'b10101; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11011; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 7,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b00110; // Expected: {'quot': 3, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 8,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 9,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b10010; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 10,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b10100; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 11,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b10101; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 12,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b00110; // Expected: {'quot': 2, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 13,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b11100; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 14,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b10000; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b10000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 15,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 16,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b11000; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b11000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 17,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b00100; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 18,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10000; Y = 5'b01111; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10000; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 19,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11111; Y = 5'b10100; // Expected: {'quot': 1, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11111; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 20,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00100; Y = 5'b00001; // Expected: {'quot': 4, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00100; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 21,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 22,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00100; Y = 5'b10101; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00100; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 23,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b10010; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 24,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b01100; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 25,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b00001; // Expected: {'quot': 9, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 26,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 9, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00100; Y = 5'b01010; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00100; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 27,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b11101; // Expected: {'quot': 0, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 28,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b10001; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 29,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00100; Y = 5'b10110; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00100; Y = 5'b10110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 30,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b01000; // Expected: {'quot': 2, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b01000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 31,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11000; Y = 5'b11010; // Expected: {'quot': 0, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11000; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 32,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b10011; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 33,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b00101; // Expected: {'quot': 4, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 34,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b00010; // Expected: {'quot': 15, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 35,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b00100; // Expected: {'quot': 3, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 36,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 37,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00101; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00101; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 38,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10000; Y = 5'b11101; // Expected: {'quot': 0, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10000; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 39,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b10000; // Expected: {'quot': 1, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b10000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 40,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b10110; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b10110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 41,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b00011; // Expected: {'quot': 3, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 42,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00011; Y = 5'b01000; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00011; Y = 5'b01000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 43,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 44,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b10110; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b10110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 45,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b00101; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 46,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b10001; // Expected: {'quot': 0, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 47,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b01011; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 48,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b01101; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 49,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b10010; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 50,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 51,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b00110; // Expected: {'quot': 4, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 52,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 53,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00100; Y = 5'b01011; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00100; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 54,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b00100; // Expected: {'quot': 4, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 55,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00011; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00011; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 56,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b01010; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 57,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b11100; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 58,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b01011; // Expected: {'quot': 2, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 59,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b01100; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 60,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b00111; // Expected: {'quot': 2, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 61,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 62,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b10010; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 63,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11111; Y = 5'b00101; // Expected: {'quot': 6, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11111; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 64,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b11001; // Expected: {'quot': 0, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 65,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b10001; // Expected: {'quot': 1, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 66,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b01011; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 67,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b11000; // Expected: {'quot': 0, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b11000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 68,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b01001; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 69,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b10001; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 70,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b10100; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 71,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b10010; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 72,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11011; Y = 5'b00100; // Expected: {'quot': 6, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11011; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 73,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b01010; // Expected: {'quot': 2, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 74,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11011; Y = 5'b01011; // Expected: {'quot': 2, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11011; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 75,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b00111; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 76,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b01001; // Expected: {'quot': 2, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 77,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b01010; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 78,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b00010; // Expected: {'quot': 7, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 79,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b11100; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 80,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b10010; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 81,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b11010; // Expected: {'quot': 1, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 82,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b01001; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 83,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b11001; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 84,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b00101; // Expected: {'quot': 6, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 85,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11000; Y = 5'b10100; // Expected: {'quot': 1, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11000; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 86,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b01100; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 87,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b00101; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 88,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00011; Y = 5'b11010; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00011; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 89,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00100; Y = 5'b11001; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00100; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 90,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 91,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b10011; // Expected: {'quot': 0, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 92,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b10111; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 93,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b00010; // Expected: {'quot': 5, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 94,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b01101; // Expected: {'quot': 1, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 95,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 96,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b00001; // Expected: {'quot': 20, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 97,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 20, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00100; Y = 5'b10110; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00100; Y = 5'b10110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 98,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b00010; // Expected: {'quot': 7, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 99,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b01010; // Expected: {'quot': 2, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 100,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11111; Y = 5'b00110; // Expected: {'quot': 5, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11111; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 101,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b01011; // Expected: {'quot': 2, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 102,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b00010; // Expected: {'quot': 6, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 103,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b01000; // Expected: {'quot': 3, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b01000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 104,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b01110; // Expected: {'quot': 1, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 105,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b10110; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b10110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 106,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b10101; // Expected: {'quot': 0, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 107,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b01110; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 108,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b10000; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b10000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 109,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b10010; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 110,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b11000; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b11000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 111,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b00001; // Expected: {'quot': 14, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 112,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b11100; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 113,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b10011; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 114,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b01010; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 115,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11111; Y = 5'b00100; // Expected: {'quot': 7, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11111; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 116,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b01001; // Expected: {'quot': 2, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 117,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b11101; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 118,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 119,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b00011; // Expected: {'quot': 7, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 120,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b01111; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 121,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b00100; // Expected: {'quot': 5, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 122,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b11010; // Expected: {'quot': 0, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 123,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b00110; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 124,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00011; Y = 5'b10111; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00011; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 125,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b10110; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b10110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 126,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b11000; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b11000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 127,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b01100; // Expected: {'quot': 1, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 128,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b01100; // Expected: {'quot': 1, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 129,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b01101; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 130,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00011; Y = 5'b10100; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00011; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 131,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b01110; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 132,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b10110; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b10110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 133,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b00111; // Expected: {'quot': 4, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 134,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00101; Y = 5'b10110; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00101; Y = 5'b10110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 135,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11111; Y = 5'b01110; // Expected: {'quot': 2, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11111; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 136,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b01100; // Expected: {'quot': 1, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 137,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 138,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00011; Y = 5'b01000; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00011; Y = 5'b01000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 139,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 140,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b00010; // Expected: {'quot': 11, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 141,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 11, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b01110; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 142,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b10000; // Expected: {'quot': 1, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b10000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 143,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b11101; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 144,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b10110; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b10110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 145,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b11101; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 146,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 147,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 148,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b01010; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 149,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 150,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b00010; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 151,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b01010; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 152,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b10011; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 153,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 154,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b11101; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 155,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b00100; // Expected: {'quot': 7, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 156,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b11000; // Expected: {'quot': 0, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b11000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 157,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b00111; // Expected: {'quot': 2, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 158,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b00101; // Expected: {'quot': 6, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 159,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b11001; // Expected: {'quot': 0, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 160,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b01111; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 161,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b10010; // Expected: {'quot': 1, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 162,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b00100; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 163,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b01110; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 164,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b11001; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 165,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b00111; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 166,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b10000; // Expected: {'quot': 1, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b10000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 167,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b00010; // Expected: {'quot': 7, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 168,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b11000; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b11000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 169,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b11010; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 170,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00101; Y = 5'b11100; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00101; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 171,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b01010; // Expected: {'quot': 2, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 172,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b01111; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 173,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11000; Y = 5'b01001; // Expected: {'quot': 2, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11000; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 174,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b11100; // Expected: {'quot': 0, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 175,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 176,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b01101; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 177,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b00001; // Expected: {'quot': 18, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 178,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 18, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b01101; // Expected: {'quot': 1, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 179,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b01100; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 180,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b01111; // Expected: {'quot': 2, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 181,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b10001; // Expected: {'quot': 1, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 182,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b10100; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 183,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b00111; // Expected: {'quot': 3, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 184,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b00001; // Expected: {'quot': 19, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 185,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 19, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 186,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b10010; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 187,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b10011; // Expected: {'quot': 1, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 188,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b00111; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 189,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00011; Y = 5'b10010; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00011; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 190,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b11001; // Expected: {'quot': 0, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 191,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00100; Y = 5'b00110; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00100; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 192,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11011; Y = 5'b01100; // Expected: {'quot': 2, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11011; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 193,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b01101; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 194,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b01111; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 195,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11011; Y = 5'b01100; // Expected: {'quot': 2, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11011; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 196,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b10111; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 197,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b10111; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 198,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b01101; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 199,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10000; Y = 5'b00111; // Expected: {'quot': 2, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10000; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 200,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 201,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 202,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b10001; // Expected: {'quot': 0, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 203,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b10101; // Expected: {'quot': 0, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 204,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10000; Y = 5'b00011; // Expected: {'quot': 5, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10000; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 205,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11000; Y = 5'b00110; // Expected: {'quot': 4, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11000; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 206,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b01011; // Expected: {'quot': 2, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 207,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b00010; // Expected: {'quot': 14, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 208,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b11001; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 209,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b01000; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b01000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 210,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b11101; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 211,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00101; Y = 5'b00101; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00101; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 212,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b10011; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 213,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11011; Y = 5'b01101; // Expected: {'quot': 2, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11011; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 214,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b10110; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b10110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 215,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b10001; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 216,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b00011; // Expected: {'quot': 3, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 217,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10000; Y = 5'b01011; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10000; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 218,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b01010; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 219,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b10101; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 220,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b10111; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 221,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00011; Y = 5'b10001; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00011; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 222,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b00101; // Expected: {'quot': 4, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 223,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10000; Y = 5'b10101; // Expected: {'quot': 0, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10000; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 224,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b11101; // Expected: {'quot': 0, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 225,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b00100; // Expected: {'quot': 2, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 226,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b00010; // Expected: {'quot': 15, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 227,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11000; Y = 5'b01100; // Expected: {'quot': 2, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11000; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 228,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b01110; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 229,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b00110; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 230,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b01010; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 231,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b11100; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 232,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b10010; // Expected: {'quot': 0, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 233,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b10000; // Expected: {'quot': 1, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b10000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 234,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b11001; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 235,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b00110; // Expected: {'quot': 3, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 236,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b01011; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 237,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 238,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b01010; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 239,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b01001; // Expected: {'quot': 2, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 240,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b00111; // Expected: {'quot': 4, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 241,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b00010; // Expected: {'quot': 8, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 242,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b10100; // Expected: {'quot': 0, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 243,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11111; Y = 5'b11100; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11111; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 244,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b10111; // Expected: {'quot': 0, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 245,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b00100; // Expected: {'quot': 3, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 246,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b10001; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 247,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b00101; // Expected: {'quot': 5, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 248,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 249,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b00001; // Expected: {'quot': 7, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 250,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b00001; // Expected: {'quot': 9, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 251,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 9, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b11000; // Expected: {'quot': 0, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b11000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 252,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11011; Y = 5'b11101; // Expected: {'quot': 0, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11011; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 253,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b01110; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 254,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b11010; // Expected: {'quot': 0, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 255,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b01101; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 256,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b11100; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 257,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b10011; // Expected: {'quot': 1, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 258,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b01001; // Expected: {'quot': 2, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 259,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b01110; // Expected: {'quot': 1, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 260,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b01111; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 261,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b10011; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 262,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00100; Y = 5'b01111; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00100; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 263,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b01011; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 264,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b10000; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b10000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 265,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11011; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11011; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 266,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11011; Y = 5'b10101; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11011; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 267,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b10011; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 268,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b01111; // Expected: {'quot': 0, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 269,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11000; Y = 5'b01100; // Expected: {'quot': 2, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11000; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 270,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 271,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b01011; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 272,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b00001; // Expected: {'quot': 28, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 273,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 28, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b11010; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 274,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11111; Y = 5'b11101; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11111; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 275,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b00101; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 276,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b11001; // Expected: {'quot': 1, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 277,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b01001; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 278,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 25}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 279,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b00010; // Expected: {'quot': 14, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 280,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b00001; // Expected: {'quot': 25, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 281,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 25, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b11000; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b11000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 282,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b00001; // Expected: {'quot': 10, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 283,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 10, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b11101; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 284,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b00111; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 285,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b01000; // Expected: {'quot': 2, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b01000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 286,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b00110; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 287,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00101; Y = 5'b00011; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00101; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 288,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b11101; // Expected: {'quot': 0, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 289,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b00101; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 290,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10000; Y = 5'b01010; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10000; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 291,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b10111; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 292,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b00110; // Expected: {'quot': 4, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 293,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b00011; // Expected: {'quot': 3, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 294,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b10111; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 295,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b11010; // Expected: {'quot': 0, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 296,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b01001; // Expected: {'quot': 2, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 297,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11000; Y = 5'b10111; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11000; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 298,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b01001; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 299,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 300,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11000; Y = 5'b10001; // Expected: {'quot': 1, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11000; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 301,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b10000; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b10000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 302,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b00110; // Expected: {'quot': 1, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 303,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10000; Y = 5'b01001; // Expected: {'quot': 1, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10000; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 304,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b01110; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 305,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 306,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00101; Y = 5'b01110; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00101; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 307,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b11101; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 308,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b00110; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 309,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 310,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b11101; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 311,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b00010; // Expected: {'quot': 7, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 312,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b11010; // Expected: {'quot': 0, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 313,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b11001; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 314,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b10001; // Expected: {'quot': 1, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 315,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00011; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00011; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 316,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b11010; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 317,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b00101; // Expected: {'quot': 5, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 318,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b01011; // Expected: {'quot': 1, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 319,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 320,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b10100; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 321,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11111; Y = 5'b10111; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11111; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 322,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b00011; // Expected: {'quot': 6, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 323,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b01001; // Expected: {'quot': 2, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 324,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b01010; // Expected: {'quot': 3, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 325,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b10000; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b10000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 326,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b01100; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 327,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b01010; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 328,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b00011; // Expected: {'quot': 7, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 329,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b00001; // Expected: {'quot': 18, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 330,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 18, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b11010; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 331,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b01010; // Expected: {'quot': 2, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 332,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b10000; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b10000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 333,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b10101; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 334,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 335,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b11100; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 336,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b01100; // Expected: {'quot': 2, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 337,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b00101; // Expected: {'quot': 4, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 338,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b00111; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 339,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b00101; // Expected: {'quot': 4, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 340,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b00001; // Expected: {'quot': 13, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 341,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b11100; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 342,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b01011; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 343,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 344,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b01110; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 345,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b01101; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 346,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b10100; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 347,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 348,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b00111; // Expected: {'quot': 2, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 349,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b10000; // Expected: {'quot': 0, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b10000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 350,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b11100; // Expected: {'quot': 0, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 351,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00011; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00011; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 352,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b10101; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 353,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b01110; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 354,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b00100; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 355,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 356,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b00111; // Expected: {'quot': 3, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 357,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b10100; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 358,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00011; Y = 5'b01001; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00011; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 359,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b00110; // Expected: {'quot': 2, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 360,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b01110; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 361,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b01101; // Expected: {'quot': 2, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 362,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b10011; // Expected: {'quot': 1, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 363,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b10100; // Expected: {'quot': 0, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 364,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00101; Y = 5'b11000; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00101; Y = 5'b11000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 365,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b00110; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 366,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00101; Y = 5'b00101; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00101; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 367,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b00100; // Expected: {'quot': 2, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 368,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b00010; // Expected: {'quot': 9, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 369,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 9, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b10010; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 370,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b11100; // Expected: {'quot': 0, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 371,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b10111; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 372,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b00001; // Expected: {'quot': 15, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 373,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b01011; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 374,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b11001; // Expected: {'quot': 0, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 375,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b10000; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b10000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 376,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b01100; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 377,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00101; Y = 5'b00110; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00101; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 378,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00011; Y = 5'b00100; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00011; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 379,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11111; Y = 5'b11000; // Expected: {'quot': 1, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11111; Y = 5'b11000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 380,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b00111; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 381,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b10100; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 382,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b10110; // Expected: {'quot': 0, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b10110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 383,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b00100; // Expected: {'quot': 3, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 384,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b01001; // Expected: {'quot': 2, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 385,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b00011; // Expected: {'quot': 6, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 386,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b11100; // Expected: {'quot': 0, 'rem': 25}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 387,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11000; Y = 5'b10011; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11000; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 388,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b00111; // Expected: {'quot': 3, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 389,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b10010; // Expected: {'quot': 0, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 390,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b00010; // Expected: {'quot': 14, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 391,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00011; Y = 5'b00101; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00011; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 392,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b00111; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 393,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b00111; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 394,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00011; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00011; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 395,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b11001; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 396,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b11101; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 397,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b01000; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b01000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 398,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 399,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b10001; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 400,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b10111; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 401,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b01101; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 402,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b01000; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b01000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 403,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b10111; // Expected: {'quot': 0, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 404,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b10111; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 405,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11011; Y = 5'b00011; // Expected: {'quot': 9, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11011; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 406,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 9, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b01011; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 407,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11011; Y = 5'b11001; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11011; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 408,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b01010; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 409,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b10101; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 410,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10000; Y = 5'b01101; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10000; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 411,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b11101; // Expected: {'quot': 0, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 412,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b00110; // Expected: {'quot': 3, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 413,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b01101; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 414,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b11101; // Expected: {'quot': 0, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 415,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b00110; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 416,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b01100; // Expected: {'quot': 2, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 417,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00011; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00011; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 418,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11111; Y = 5'b10011; // Expected: {'quot': 1, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11111; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 419,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b00100; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 420,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b01101; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 421,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b01110; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 422,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 423,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b11010; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 424,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 425,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00011; Y = 5'b10001; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00011; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 426,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00100; Y = 5'b00111; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00100; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 427,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b10011; // Expected: {'quot': 0, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 428,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b00110; // Expected: {'quot': 3, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 429,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b01001; // Expected: {'quot': 1, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 430,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00101; Y = 5'b01111; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00101; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 431,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 432,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b10000; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b10000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 433,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 434,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 435,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b00001; // Expected: {'quot': 15, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 436,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b11101; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 437,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00100; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00100; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 438,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00100; Y = 5'b10011; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00100; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 439,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 25}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 440,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b10000; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b10000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 441,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 442,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b01111; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 443,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b10001; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 444,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b00011; // Expected: {'quot': 6, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 445,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b01111; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 446,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b10001; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 447,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b11000; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b11000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 448,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b10111; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 449,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b01100; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 450,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b01001; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 451,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11111; Y = 5'b00001; // Expected: {'quot': 31, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11111; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 452,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 31, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b01000; // Expected: {'quot': 2, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b01000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 453,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b01011; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 454,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b11001; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 455,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b00011; // Expected: {'quot': 4, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 456,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b01010; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 457,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b00010; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 458,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 459,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b01110; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 460,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b10111; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 461,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b10010; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 462,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b10011; // Expected: {'quot': 0, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 463,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00011; Y = 5'b01000; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00011; Y = 5'b01000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 464,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b00001; // Expected: {'quot': 21, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 465,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 21, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b01101; // Expected: {'quot': 2, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 466,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b11001; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 467,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b00111; // Expected: {'quot': 3, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 468,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b00111; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 469,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b10010; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 470,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 471,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 472,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b00101; // Expected: {'quot': 4, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 473,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b10100; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 474,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11000; Y = 5'b10110; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11000; Y = 5'b10110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 475,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b01011; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 476,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10000; Y = 5'b01010; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10000; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 477,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00101; Y = 5'b01011; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00101; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 478,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b10101; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 479,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 480,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b01110; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 481,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b00100; // Expected: {'quot': 3, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 482,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b10010; // Expected: {'quot': 1, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 483,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b11001; // Expected: {'quot': 0, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 484,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11000; Y = 5'b10011; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11000; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 485,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 486,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b10001; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 487,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11111; Y = 5'b11010; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11111; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 488,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b00100; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 489,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b00001; // Expected: {'quot': 7, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 490,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b10011; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 491,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b11000; // Expected: {'quot': 0, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b11000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 492,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b00111; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 493,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b11001; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 494,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 495,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b11010; // Expected: {'quot': 0, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 496,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b10100; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 497,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b00010; // Expected: {'quot': 6, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 498,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 499,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b00011; // Expected: {'quot': 2, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 500,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00100; Y = 5'b11100; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00100; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 501,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b01000; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b01000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 502,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 503,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b00100; // Expected: {'quot': 7, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 504,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b00100; // Expected: {'quot': 4, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 505,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b01100; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 506,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b11100; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 507,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b01001; // Expected: {'quot': 2, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 508,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b00001; // Expected: {'quot': 22, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 509,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 22, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b10010; // Expected: {'quot': 1, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 510,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b01000; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b01000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 511,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b00001; // Expected: {'quot': 7, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 512,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b11101; // Expected: {'quot': 0, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 513,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b00100; // Expected: {'quot': 4, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 514,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b10111; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 515,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00011; Y = 5'b01010; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00011; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 516,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b10100; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 517,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b01001; // Expected: {'quot': 1, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 518,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b11100; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 519,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b01010; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 520,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b10101; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 521,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b10111; // Expected: {'quot': 0, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 522,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b10100; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 523,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b10011; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 524,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b00011; // Expected: {'quot': 2, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 525,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b01011; // Expected: {'quot': 2, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 526,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b00100; // Expected: {'quot': 2, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 527,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b00010; // Expected: {'quot': 15, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 528,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b10110; // Expected: {'quot': 0, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b10110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 529,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b11001; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 530,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b10101; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 531,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11111; Y = 5'b00011; // Expected: {'quot': 10, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11111; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 532,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b01000; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b01000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 533,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b10100; // Expected: {'quot': 1, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 534,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b01010; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 535,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b01101; // Expected: {'quot': 1, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 536,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11111; Y = 5'b00110; // Expected: {'quot': 5, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11111; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 537,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b00011; // Expected: {'quot': 6, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 538,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b11001; // Expected: {'quot': 0, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 539,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b01110; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 540,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 541,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11111; Y = 5'b11011; // Expected: {'quot': 1, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11111; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 542,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b00001; // Expected: {'quot': 26, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 543,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 26, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b01000; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b01000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 544,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b00010; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 545,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b01101; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 546,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 547,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11000; Y = 5'b11100; // Expected: {'quot': 0, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11000; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 548,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b10010; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 549,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b00001; // Expected: {'quot': 25, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 550,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 25, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10000; Y = 5'b10111; // Expected: {'quot': 0, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10000; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 551,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b01011; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 552,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10000; Y = 5'b11001; // Expected: {'quot': 0, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10000; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 553,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b01010; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 554,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b10001; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 555,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b01101; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 556,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10000; Y = 5'b10101; // Expected: {'quot': 0, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10000; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 557,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b10100; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 558,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b01110; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 559,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b01110; // Expected: {'quot': 1, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 560,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11011; Y = 5'b01010; // Expected: {'quot': 2, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11011; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 561,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00011; Y = 5'b10000; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00011; Y = 5'b10000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 562,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b11000; // Expected: {'quot': 0, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b11000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 563,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b01010; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 564,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10000; Y = 5'b10111; // Expected: {'quot': 0, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10000; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 565,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b01001; // Expected: {'quot': 2, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 566,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00100; Y = 5'b00011; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00100; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 567,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b00101; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 568,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b01011; // Expected: {'quot': 2, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 569,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11011; Y = 5'b01110; // Expected: {'quot': 1, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11011; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 570,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00101; Y = 5'b10100; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00101; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 571,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b00110; // Expected: {'quot': 4, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 572,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b01010; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 573,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b00110; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 574,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b00001; // Expected: {'quot': 28, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 575,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 28, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00101; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00101; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 576,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b01111; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 577,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 578,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b11101; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 579,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b10110; // Expected: {'quot': 0, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b10110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 580,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b01011; // Expected: {'quot': 1, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 581,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11000; Y = 5'b11000; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11000; Y = 5'b11000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 582,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b01101; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 583,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b01110; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 584,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00100; Y = 5'b11010; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00100; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 585,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b10110; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b10110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 586,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10000; Y = 5'b00110; // Expected: {'quot': 2, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10000; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 587,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b11101; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 588,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b01000; // Expected: {'quot': 3, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b01000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 589,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 25}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 590,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b01101; // Expected: {'quot': 1, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 591,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b01111; // Expected: {'quot': 2, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 592,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b00111; // Expected: {'quot': 4, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 593,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b10110; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b10110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 594,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b01001; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 595,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b11001; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 596,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b01010; // Expected: {'quot': 2, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 597,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b11001; // Expected: {'quot': 0, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 598,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b10011; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 599,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b00110; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 600,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b11010; // Expected: {'quot': 0, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 601,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b10011; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 602,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b10110; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b10110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 603,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10000; Y = 5'b01111; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10000; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 604,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b01010; // Expected: {'quot': 2, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 605,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11000; Y = 5'b00111; // Expected: {'quot': 3, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11000; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 606,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b11001; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 607,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11011; Y = 5'b00111; // Expected: {'quot': 3, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11011; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 608,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b10100; // Expected: {'quot': 1, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 609,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b10001; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 610,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b01011; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 611,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b00100; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 612,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b00011; // Expected: {'quot': 5, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 613,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10000; Y = 5'b10100; // Expected: {'quot': 0, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10000; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 614,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11011; Y = 5'b10111; // Expected: {'quot': 1, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11011; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 615,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00101; Y = 5'b10101; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00101; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 616,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b10100; // Expected: {'quot': 1, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 617,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b10100; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 618,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11111; Y = 5'b10101; // Expected: {'quot': 1, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11111; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 619,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11000; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11000; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 620,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b01100; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 621,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b10101; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 622,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10000; Y = 5'b10100; // Expected: {'quot': 0, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10000; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 623,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11011; Y = 5'b01001; // Expected: {'quot': 3, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11011; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 624,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b10110; // Expected: {'quot': 0, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b10110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 625,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b00010; // Expected: {'quot': 7, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 626,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11011; Y = 5'b01111; // Expected: {'quot': 1, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11011; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 627,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b10100; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 628,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b11110; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 629,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b01101; // Expected: {'quot': 1, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 630,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b11100; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 631,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b10001; // Expected: {'quot': 1, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 632,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b01100; // Expected: {'quot': 1, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 633,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b11010; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 634,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b01011; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 635,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b10011; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 636,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b01100; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 637,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b11000; // Expected: {'quot': 0, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b11000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 638,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b10101; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 639,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11000; Y = 5'b10001; // Expected: {'quot': 1, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11000; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 640,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b10100; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 641,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b10011; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 642,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00101; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00101; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 643,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b00010; // Expected: {'quot': 14, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 644,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b00001; // Expected: {'quot': 15, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 645,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b01011; // Expected: {'quot': 2, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 646,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 647,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b10100; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 648,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 649,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b01011; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 650,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b01011; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 651,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b00001; // Expected: {'quot': 30, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 652,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 30, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b10101; // Expected: {'quot': 0, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 653,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b11101; // Expected: {'quot': 0, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 654,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b11101; // Expected: {'quot': 0, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 655,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b11000; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b11000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 656,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11000; Y = 5'b01100; // Expected: {'quot': 2, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11000; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 657,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b10100; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 658,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b10001; // Expected: {'quot': 0, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 659,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11011; Y = 5'b11100; // Expected: {'quot': 0, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11011; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 660,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b00101; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 661,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b01100; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 662,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b01011; // Expected: {'quot': 2, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 663,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b11001; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 664,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b00111; // Expected: {'quot': 4, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 665,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00100; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00100; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 666,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b01000; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b01000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 667,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b00100; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 668,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b01101; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 669,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b11100; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 670,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b10111; // Expected: {'quot': 1, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 671,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b00101; // Expected: {'quot': 1, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 672,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b01010; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 673,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b11010; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 674,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b00110; // Expected: {'quot': 2, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 675,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b10101; // Expected: {'quot': 0, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 676,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b11001; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 677,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b01111; // Expected: {'quot': 1, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 678,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b11010; // Expected: {'quot': 0, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 679,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b01011; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 680,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b11001; // Expected: {'quot': 0, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 681,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b10000; // Expected: {'quot': 1, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b10000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 682,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b11010; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 683,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b00010; // Expected: {'quot': 8, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 684,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00101; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00101; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 685,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b01110; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 686,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b10011; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 687,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b01010; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 688,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10000; Y = 5'b00101; // Expected: {'quot': 3, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10000; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 689,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b01110; // Expected: {'quot': 2, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 690,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 25}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 691,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b01011; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 692,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b01000; // Expected: {'quot': 2, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b01000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 693,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 694,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b10101; // Expected: {'quot': 0, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 695,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 696,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10000; Y = 5'b00100; // Expected: {'quot': 4, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10000; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 697,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b00011; // Expected: {'quot': 2, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 698,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11000; Y = 5'b00100; // Expected: {'quot': 6, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11000; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 699,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b10111; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 700,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b10010; // Expected: {'quot': 1, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 701,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b10011; // Expected: {'quot': 0, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 702,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b10001; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 703,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b00101; // Expected: {'quot': 1, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 704,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b11010; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 705,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b10010; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 706,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b11000; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b11000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 707,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b01011; // Expected: {'quot': 1, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 708,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11111; Y = 5'b01001; // Expected: {'quot': 3, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11111; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 709,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11000; Y = 5'b11101; // Expected: {'quot': 0, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11000; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 710,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b10101; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 711,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11000; Y = 5'b10011; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11000; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 712,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b11001; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 713,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b00110; // Expected: {'quot': 4, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 714,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b10001; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 715,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b11000; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b11000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 716,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b10100; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 717,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b00010; // Expected: {'quot': 4, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 718,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b01111; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 719,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00100; Y = 5'b10000; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00100; Y = 5'b10000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 720,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b00010; // Expected: {'quot': 9, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 721,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 9, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10000; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10000; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 722,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b01001; // Expected: {'quot': 2, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 723,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b00001; // Expected: {'quot': 23, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 724,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 23, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b01101; // Expected: {'quot': 2, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 725,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 726,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b10101; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 727,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00011; Y = 5'b00100; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00011; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 728,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10000; Y = 5'b11100; // Expected: {'quot': 0, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10000; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 729,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b01010; // Expected: {'quot': 1, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 730,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00101; Y = 5'b01000; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00101; Y = 5'b01000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 731,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b01110; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 732,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b10011; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 733,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b11011; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 734,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b01010; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 735,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b00001; // Expected: {'quot': 26, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 736,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 26, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b10111; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 737,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b00011; // Expected: {'quot': 6, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 738,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00011; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00011; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 739,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 740,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b11000; // Expected: {'quot': 0, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b11000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 741,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b10100; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 742,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b00100; // Expected: {'quot': 4, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 743,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b10001; // Expected: {'quot': 1, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 744,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11111; Y = 5'b00101; // Expected: {'quot': 6, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11111; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 745,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b00011; // Expected: {'quot': 4, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 746,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b00110; // Expected: {'quot': 2, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 747,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b01000; // Expected: {'quot': 3, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b01000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 748,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b11100; // Expected: {'quot': 0, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 749,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00011; Y = 5'b01010; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00011; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 750,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b10111; // Expected: {'quot': 0, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 751,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b00101; // Expected: {'quot': 2, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 752,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11000; Y = 5'b11101; // Expected: {'quot': 0, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11000; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 753,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00101; Y = 5'b01101; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00101; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 754,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 755,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b00101; // Expected: {'quot': 3, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 756,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b00001; // Expected: {'quot': 23, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 757,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 23, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b00001; // Expected: {'quot': 22, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 758,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 22, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00100; Y = 5'b01010; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00100; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 759,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11011; Y = 5'b01010; // Expected: {'quot': 2, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11011; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 760,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b10110; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b10110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 761,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 762,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11000; Y = 5'b00001; // Expected: {'quot': 24, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11000; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 763,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 24, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b11011; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 764,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b01110; // Expected: {'quot': 1, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 765,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b11000; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b11000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 766,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b11101; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 767,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00100; Y = 5'b10101; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00100; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 768,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b10110; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b10110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 769,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b01010; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 770,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b01101; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 771,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b10001; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 772,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 773,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b10100; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 774,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00100; Y = 5'b11010; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00100; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 775,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b10011; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 776,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b11101; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 777,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b01110; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 778,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 779,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11000; Y = 5'b00111; // Expected: {'quot': 3, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11000; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 780,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b10010; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 781,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b10100; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 782,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b11010; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 783,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b01110; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 784,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11011; Y = 5'b00110; // Expected: {'quot': 4, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11011; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 785,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b01001; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 786,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00101; Y = 5'b11101; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00101; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 787,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b10010; // Expected: {'quot': 0, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 788,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b11000; // Expected: {'quot': 0, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b11000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 789,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11111; Y = 5'b01000; // Expected: {'quot': 3, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11111; Y = 5'b01000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 790,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b10010; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 791,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 792,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b10011; // Expected: {'quot': 0, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 793,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11111; Y = 5'b11010; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11111; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 794,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b01000; // Expected: {'quot': 2, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b01000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 795,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b10111; // Expected: {'quot': 1, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 796,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b01111; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 797,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b10111; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 798,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b10010; // Expected: {'quot': 1, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 799,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b10111; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 800,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b00011; // Expected: {'quot': 8, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 801,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00101; Y = 5'b01110; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00101; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 802,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b01100; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 803,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00101; Y = 5'b00110; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00101; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 804,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b11100; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 805,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b00010; // Expected: {'quot': 14, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 806,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b11010; // Expected: {'quot': 0, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 807,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b10010; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 808,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b11010; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 809,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00101; Y = 5'b10110; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00101; Y = 5'b10110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 810,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11011; Y = 5'b11100; // Expected: {'quot': 0, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11011; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 811,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b10000; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b10000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 812,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b11010; // Expected: {'quot': 0, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 813,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b00110; // Expected: {'quot': 4, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 814,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b00100; // Expected: {'quot': 5, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 815,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b10000; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b10000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 816,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11011; Y = 5'b00110; // Expected: {'quot': 4, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11011; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 817,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b00101; // Expected: {'quot': 4, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 818,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b01110; // Expected: {'quot': 2, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 819,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b11100; // Expected: {'quot': 0, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 820,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b00111; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 821,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11011; Y = 5'b11010; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11011; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 822,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b00100; // Expected: {'quot': 3, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 823,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b10011; // Expected: {'quot': 1, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 824,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b01110; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 825,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b11010; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 826,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 827,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b10110; // Expected: {'quot': 1, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b10110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 828,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b01010; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 829,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b00111; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 830,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b01100; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 831,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b01000; // Expected: {'quot': 3, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b01000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 832,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00100; Y = 5'b10011; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00100; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 833,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b01100; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 834,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b01001; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 835,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b01011; // Expected: {'quot': 2, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 836,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b01010; // Expected: {'quot': 2, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 837,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b11010; // Expected: {'quot': 1, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 838,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b10100; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 839,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 840,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b00001; // Expected: {'quot': 19, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 841,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 19, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11000; Y = 5'b00101; // Expected: {'quot': 4, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11000; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 842,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b11000; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b11000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 843,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b11101; // Expected: {'quot': 0, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 844,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b00111; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 845,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b10000; // Expected: {'quot': 1, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b10000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 846,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b01101; // Expected: {'quot': 1, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 847,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b10101; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 848,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b00110; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 849,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 850,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b01111; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 851,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b00101; // Expected: {'quot': 3, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 852,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b01100; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 853,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b00001; // Expected: {'quot': 22, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 854,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 22, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b11100; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 855,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11111; Y = 5'b10000; // Expected: {'quot': 1, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11111; Y = 5'b10000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 856,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10011; Y = 5'b00011; // Expected: {'quot': 6, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10011; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 857,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b00011; // Expected: {'quot': 4, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 858,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00011; Y = 5'b00111; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00011; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 859,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11111; Y = 5'b01100; // Expected: {'quot': 2, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11111; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 860,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b01111; // Expected: {'quot': 1, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 861,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b00110; // Expected: {'quot': 2, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 862,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b01010; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 863,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b10011; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 864,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b10001; // Expected: {'quot': 0, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 865,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b01100; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 866,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00101; Y = 5'b10101; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00101; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 867,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b00010; // Expected: {'quot': 11, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 868,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 11, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b10101; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 869,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 870,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b01101; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 871,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11011; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11011; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 872,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b00110; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 873,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b00011; // Expected: {'quot': 2, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 874,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b01010; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 875,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b10100; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b10100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 876,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b10000; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b10000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 877,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b00010; // Expected: {'quot': 10, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 878,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b10101; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 879,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b00100; // Expected: {'quot': 7, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 880,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11000; Y = 5'b10001; // Expected: {'quot': 1, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11000; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 881,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00011; Y = 5'b10110; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00011; Y = 5'b10110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 882,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b00101; // Expected: {'quot': 3, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 883,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b01000; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b01000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 884,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01110; Y = 5'b00111; // Expected: {'quot': 2, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01110; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 885,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 886,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b00101; // Expected: {'quot': 2, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 887,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b01001; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 888,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b10001; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 889,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b01101; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 890,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b01101; // Expected: {'quot': 1, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 891,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10000; Y = 5'b11001; // Expected: {'quot': 0, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10000; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 892,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b01101; // Expected: {'quot': 2, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 893,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b01111; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 894,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11111; Y = 5'b01110; // Expected: {'quot': 2, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11111; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 895,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b11010; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b11010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 896,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b00110; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 897,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b10010; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 898,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b00100; // Expected: {'quot': 5, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 899,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b10101; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 900,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b01110; // Expected: {'quot': 1, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 901,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b10101; // Expected: {'quot': 1, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 902,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11011; Y = 5'b01110; // Expected: {'quot': 1, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11011; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 903,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b00011; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 904,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b10010; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 905,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b01111; // Expected: {'quot': 1, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 906,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b01001; // Expected: {'quot': 3, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 907,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b01111; // Expected: {'quot': 1, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 908,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b01001; // Expected: {'quot': 3, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b01001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 909,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b00001; // Expected: {'quot': 2, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 910,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b11000; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b11000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 911,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b11101; // Expected: {'quot': 0, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 912,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b11110; // Expected: {'quot': 0, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b11110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 913,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b01111; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 914,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b01111; // Expected: {'quot': 1, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 915,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b10110; // Expected: {'quot': 0, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b10110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 916,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11000; Y = 5'b01101; // Expected: {'quot': 1, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11000; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 917,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10000; Y = 5'b10101; // Expected: {'quot': 0, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10000; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 918,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11111; Y = 5'b10001; // Expected: {'quot': 1, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11111; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 919,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b00010; // Expected: {'quot': 14, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 920,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b11000; // Expected: {'quot': 0, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b11000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 921,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b10001; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 922,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b11100; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 923,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b11001; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 924,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b01101; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 925,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b11001; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 926,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b00100; // Expected: {'quot': 2, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 927,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b10000; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b10000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 928,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b11100; // Expected: {'quot': 0, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 929,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b10011; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 930,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b00110; // Expected: {'quot': 3, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 931,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b00011; // Expected: {'quot': 8, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 932,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00100; Y = 5'b00010; // Expected: {'quot': 2, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00100; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 933,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b01111; // Expected: {'quot': 1, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 934,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11000; Y = 5'b01101; // Expected: {'quot': 1, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11000; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 935,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b01100; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 936,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b00010; // Expected: {'quot': 12, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 937,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b11100; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 938,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b00001; // Expected: {'quot': 12, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 939,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 12, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b00011; // Expected: {'quot': 5, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b00011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 940,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00110; Y = 5'b01101; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00110; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 941,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b01100; // Expected: {'quot': 2, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 942,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b00100; // Expected: {'quot': 7, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 943,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b10010; // Expected: {'quot': 0, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 944,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 945,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b01011; // Expected: {'quot': 2, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b01011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 946,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b10101; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 947,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00100; Y = 5'b01010; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00100; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 948,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b10011; // Expected: {'quot': 1, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 949,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00100; Y = 5'b10101; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00100; Y = 5'b10101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 950,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b11001; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 951,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10101; Y = 5'b10011; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10101; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 952,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b10001; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 953,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b01010; // Expected: {'quot': 3, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 954,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b01100; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 955,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b01010; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 956,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11101; Y = 5'b11101; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11101; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 957,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00001; Y = 5'b00010; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00001; Y = 5'b00010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 958,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00000; Y = 5'b11000; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00000; Y = 5'b11000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 959,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b01010; // Expected: {'quot': 2, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 960,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10111; Y = 5'b10111; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10111; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 961,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11010; Y = 5'b11100; // Expected: {'quot': 0, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11010; Y = 5'b11100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 962,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00010; Y = 5'b00101; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00010; Y = 5'b00101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 963,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00011; Y = 5'b10000; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00011; Y = 5'b10000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 964,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b11101; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 965,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b10000; // Expected: {'quot': 1, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b10000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 966,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01001; Y = 5'b01000; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01001; Y = 5'b01000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 967,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b10001; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 968,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00101; Y = 5'b01101; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00101; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 969,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01010; Y = 5'b10001; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01010; Y = 5'b10001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 970,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10010; Y = 5'b00110; // Expected: {'quot': 3, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10010; Y = 5'b00110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 971,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b00111; // Expected: {'quot': 3, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b00111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 972,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11111; Y = 5'b10011; // Expected: {'quot': 1, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11111; Y = 5'b10011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 973,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10001; Y = 5'b11001; // Expected: {'quot': 0, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10001; Y = 5'b11001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 974,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10100; Y = 5'b01100; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10100; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 975,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b01110; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 976,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01111; Y = 5'b10010; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01111; Y = 5'b10010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 977,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b10110; Y = 5'b11101; // Expected: {'quot': 0, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b10110; Y = 5'b11101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 978,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b01101; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b01101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 979,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00011; Y = 5'b01110; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00011; Y = 5'b01110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 980,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b10111; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b10111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 981,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11001; Y = 5'b00001; // Expected: {'quot': 25, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11001; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 982,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 25, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01101; Y = 5'b00001; // Expected: {'quot': 13, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01101; Y = 5'b00001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 983,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11011; Y = 5'b10000; // Expected: {'quot': 1, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11011; Y = 5'b10000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 984,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b01100; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b01100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 985,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01000; Y = 5'b01111; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01000; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 986,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b00111; Y = 5'b01010; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b00111; Y = 5'b01010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 987,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11110; Y = 5'b11111; // Expected: {'quot': 0, 'rem': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11110; Y = 5'b11111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 988,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01011; Y = 5'b00100; // Expected: {'quot': 2, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01011; Y = 5'b00100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 989,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b01100; Y = 5'b11011; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b01100; Y = 5'b11011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 990,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 5'b11100; Y = 5'b01111; // Expected: {'quot': 1, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 5'b11100; Y = 5'b01111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 991,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        $finish;
    end
  
endmodule