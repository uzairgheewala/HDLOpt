
`timescale 1ns / 1ps

module tb_N8_carry_select_adder;

    // Parameters
    
    parameter N = 8;
    
     
    // Inputs
    
    reg  [7:0] a;
    
    reg  [7:0] b;
    
    reg   cin;
    
    
    // Outputs
    
    wire  [7:0] sum;
    
    wire   cout;
    
    
    // Instantiate the Unit Under Test (UUT)
    carry_select_adder  #( N ) uut (
        
        .a(a),
        
        .b(b),
        
        .cin(cin),
        
        
        .sum(sum),
        
        .cout(cout)
        
    );
    
    initial begin
        // Initialize Inputs
        
        a = 0;
        
        b = 0;
        
        cin = 0;
        
    
        // Wait for global reset
        #100;
    
        // Stimuli
        
        a = 8'b00010011; b = 8'b00111001; cin = 1'b0; // Expected: {'sum': 76, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b00111001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 0,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 76, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010100; b = 8'b10100000; cin = 1'b0; // Expected: {'sum': 52, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010100; b = 8'b10100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 52, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011100; b = 8'b10011110; cin = 1'b0; // Expected: {'sum': 122, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011100; b = 8'b10011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 122, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100010; b = 8'b10111111; cin = 1'b0; // Expected: {'sum': 97, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100010; b = 8'b10111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 97, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110000; b = 8'b10110000; cin = 1'b1; // Expected: {'sum': 225, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110000; b = 8'b10110000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 4,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 225, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b00000000; cin = 1'b0; // Expected: {'sum': 228, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b00000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 5,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 228, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b11110000; cin = 1'b1; // Expected: {'sum': 167, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b11110000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 6,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 167, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b11000111; cin = 1'b0; // Expected: {'sum': 118, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b11000111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 7,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 118, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b10101010; cin = 1'b0; // Expected: {'sum': 36, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b10101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 8,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 36, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b11100000; cin = 1'b1; // Expected: {'sum': 254, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b11100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 9,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 254, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100111; b = 8'b11010101; cin = 1'b1; // Expected: {'sum': 61, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100111; b = 8'b11010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 10,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 61, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001000; b = 8'b11000100; cin = 1'b0; // Expected: {'sum': 140, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001000; b = 8'b11000100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 11,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 140, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111101; b = 8'b01010000; cin = 1'b1; // Expected: {'sum': 78, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111101; b = 8'b01010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 12,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 78, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100001; b = 8'b01010001; cin = 1'b1; // Expected: {'sum': 115, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100001; b = 8'b01010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 13,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 115, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001001; b = 8'b01101100; cin = 1'b0; // Expected: {'sum': 53, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001001; b = 8'b01101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 14,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 53, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011101; b = 8'b10110011; cin = 1'b1; // Expected: {'sum': 145, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011101; b = 8'b10110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 15,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 145, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b01001010; cin = 1'b0; // Expected: {'sum': 76, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b01001010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 16,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 76, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b00000011; cin = 1'b1; // Expected: {'sum': 223, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b00000011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 17,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 223, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111000; b = 8'b00101100; cin = 1'b0; // Expected: {'sum': 36, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111000; b = 8'b00101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 18,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 36, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b01100111; cin = 1'b1; // Expected: {'sum': 73, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b01100111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 19,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 73, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b01000001; cin = 1'b1; // Expected: {'sum': 172, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b01000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 20,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 172, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b11100101; cin = 1'b1; // Expected: {'sum': 19, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b11100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 21,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 19, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b10000010; cin = 1'b0; // Expected: {'sum': 58, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b10000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 22,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 58, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001011; b = 8'b01101111; cin = 1'b0; // Expected: {'sum': 122, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001011; b = 8'b01101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 23,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 122, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b10110001; cin = 1'b1; // Expected: {'sum': 166, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b10110001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 24,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 166, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b00111011; cin = 1'b0; // Expected: {'sum': 58, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b00111011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 25,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 58, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b01110110; cin = 1'b0; // Expected: {'sum': 48, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b01110110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 26,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 48, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b01010110; cin = 1'b0; // Expected: {'sum': 241, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b01010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 27,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 241, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111110; b = 8'b00100110; cin = 1'b1; // Expected: {'sum': 101, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111110; b = 8'b00100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 28,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 101, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b01101001; cin = 1'b1; // Expected: {'sum': 240, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b01101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 29,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 240, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100110; b = 8'b01011001; cin = 1'b1; // Expected: {'sum': 128, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100110; b = 8'b01011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 30,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 128, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011100; b = 8'b01111100; cin = 1'b1; // Expected: {'sum': 89, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011100; b = 8'b01111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 31,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 89, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011010; b = 8'b00010011; cin = 1'b0; // Expected: {'sum': 109, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011010; b = 8'b00010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 32,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 109, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b11011001; cin = 1'b0; // Expected: {'sum': 225, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b11011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 33,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 225, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b11110000; cin = 1'b0; // Expected: {'sum': 38, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b11110000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 34,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 38, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b10111110; cin = 1'b1; // Expected: {'sum': 232, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b10111110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 35,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 232, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011001; b = 8'b00110000; cin = 1'b0; // Expected: {'sum': 137, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011001; b = 8'b00110000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 36,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 137, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011010; b = 8'b01000011; cin = 1'b1; // Expected: {'sum': 30, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011010; b = 8'b01000011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 37,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 30, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b00100011; cin = 1'b0; // Expected: {'sum': 52, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b00100011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 38,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 52, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b00011011; cin = 1'b1; // Expected: {'sum': 194, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b00011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 39,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 194, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b01111010; cin = 1'b1; // Expected: {'sum': 248, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b01111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 40,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 248, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b10000000; cin = 1'b1; // Expected: {'sum': 251, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b10000000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 41,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 251, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111000; b = 8'b10101001; cin = 1'b0; // Expected: {'sum': 161, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111000; b = 8'b10101001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 42,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 161, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b10011000; cin = 1'b0; // Expected: {'sum': 162, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b10011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 43,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 162, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b00001101; cin = 1'b0; // Expected: {'sum': 241, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b00001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 44,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 241, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101111; b = 8'b01001110; cin = 1'b1; // Expected: {'sum': 190, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101111; b = 8'b01001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 45,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 190, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000101; b = 8'b11001010; cin = 1'b1; // Expected: {'sum': 80, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000101; b = 8'b11001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 46,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 80, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b00010000; cin = 1'b0; // Expected: {'sum': 251, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b00010000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 47,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 251, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b10011000; cin = 1'b0; // Expected: {'sum': 251, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b10011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 48,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 251, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b11100011; cin = 1'b1; // Expected: {'sum': 189, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b11100011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 49,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 189, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111101; b = 8'b00000011; cin = 1'b0; // Expected: {'sum': 0, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111101; b = 8'b00000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 50,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b10111100; cin = 1'b0; // Expected: {'sum': 187, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b10111100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 51,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 187, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101111; b = 8'b10010011; cin = 1'b1; // Expected: {'sum': 195, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101111; b = 8'b10010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 52,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 195, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b01010101; cin = 1'b1; // Expected: {'sum': 93, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b01010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 53,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 93, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010010; b = 8'b10000000; cin = 1'b0; // Expected: {'sum': 146, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010010; b = 8'b10000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 54,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 146, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b01011000; cin = 1'b1; // Expected: {'sum': 8, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b01011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 55,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 8, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b01100000; cin = 1'b1; // Expected: {'sum': 195, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b01100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 56,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 195, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001100; b = 8'b11011001; cin = 1'b0; // Expected: {'sum': 165, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001100; b = 8'b11011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 57,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 165, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b00110100; cin = 1'b0; // Expected: {'sum': 9, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b00110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 58,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 9, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100010; b = 8'b11100101; cin = 1'b1; // Expected: {'sum': 200, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100010; b = 8'b11100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 59,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 200, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b10011011; cin = 1'b0; // Expected: {'sum': 0, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b10011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 60,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b01101111; cin = 1'b0; // Expected: {'sum': 106, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b01101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 61,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 106, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110000; b = 8'b00000010; cin = 1'b0; // Expected: {'sum': 50, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110000; b = 8'b00000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 62,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 50, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b10100110; cin = 1'b0; // Expected: {'sum': 47, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b10100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 63,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 47, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b01100110; cin = 1'b1; // Expected: {'sum': 87, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b01100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 64,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 87, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101101; b = 8'b11101100; cin = 1'b0; // Expected: {'sum': 153, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101101; b = 8'b11101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 65,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 153, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001011; b = 8'b01000101; cin = 1'b1; // Expected: {'sum': 81, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001011; b = 8'b01000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 66,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 81, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001100; b = 8'b01001011; cin = 1'b0; // Expected: {'sum': 215, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001100; b = 8'b01001011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 67,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 215, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b10000111; cin = 1'b1; // Expected: {'sum': 24, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b10000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 68,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 24, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010011; b = 8'b10100000; cin = 1'b0; // Expected: {'sum': 51, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010011; b = 8'b10100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 69,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 51, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b10000111; cin = 1'b1; // Expected: {'sum': 242, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b10000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 70,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 242, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b11111000; cin = 1'b1; // Expected: {'sum': 189, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b11111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 71,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 189, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b00011001; cin = 1'b1; // Expected: {'sum': 130, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b00011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 72,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 130, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101111; b = 8'b10110101; cin = 1'b0; // Expected: {'sum': 36, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101111; b = 8'b10110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 73,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 36, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b10111000; cin = 1'b1; // Expected: {'sum': 245, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b10111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 74,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 245, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b00100110; cin = 1'b0; // Expected: {'sum': 174, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b00100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 75,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 174, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001101; b = 8'b10111111; cin = 1'b0; // Expected: {'sum': 140, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001101; b = 8'b10111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 76,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 140, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100000; b = 8'b00111110; cin = 1'b1; // Expected: {'sum': 159, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100000; b = 8'b00111110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 77,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 159, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b11101100; cin = 1'b0; // Expected: {'sum': 129, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b11101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 78,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 129, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101010; b = 8'b01100101; cin = 1'b1; // Expected: {'sum': 144, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101010; b = 8'b01100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 79,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 144, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b10110101; cin = 1'b0; // Expected: {'sum': 61, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b10110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 80,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 61, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b11011110; cin = 1'b0; // Expected: {'sum': 244, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b11011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 81,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 244, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b01010001; cin = 1'b0; // Expected: {'sum': 50, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b01010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 82,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 50, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110000; b = 8'b11011110; cin = 1'b1; // Expected: {'sum': 79, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110000; b = 8'b11011110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 83,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 79, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b01100010; cin = 1'b0; // Expected: {'sum': 58, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b01100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 84,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 58, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011001; b = 8'b00001101; cin = 1'b0; // Expected: {'sum': 166, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011001; b = 8'b00001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 85,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 166, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b01011011; cin = 1'b0; // Expected: {'sum': 121, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b01011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 86,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 121, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b00100010; cin = 1'b1; // Expected: {'sum': 155, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b00100010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 87,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 155, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100110; b = 8'b00001100; cin = 1'b1; // Expected: {'sum': 51, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100110; b = 8'b00001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 88,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 51, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b00111101; cin = 1'b1; // Expected: {'sum': 29, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b00111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 89,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 29, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001110; b = 8'b11011000; cin = 1'b0; // Expected: {'sum': 230, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001110; b = 8'b11011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 90,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 230, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b00110010; cin = 1'b0; // Expected: {'sum': 184, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b00110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 91,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 184, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b01000110; cin = 1'b0; // Expected: {'sum': 101, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b01000110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 92,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 101, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b11111011; cin = 1'b0; // Expected: {'sum': 220, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b11111011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 93,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 220, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b11000100; cin = 1'b1; // Expected: {'sum': 202, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b11000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 94,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 202, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010001; b = 8'b01011010; cin = 1'b0; // Expected: {'sum': 43, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010001; b = 8'b01011010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 95,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 43, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111111; b = 8'b10010101; cin = 1'b1; // Expected: {'sum': 213, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111111; b = 8'b10010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 96,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 213, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b01110001; cin = 1'b0; // Expected: {'sum': 120, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b01110001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 97,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 120, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b00101000; cin = 1'b1; // Expected: {'sum': 95, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b00101000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 98,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 95, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101011; b = 8'b01101001; cin = 1'b1; // Expected: {'sum': 149, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101011; b = 8'b01101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 99,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 149, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011000; b = 8'b01111010; cin = 1'b1; // Expected: {'sum': 211, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011000; b = 8'b01111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 100,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 211, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b00011001; cin = 1'b1; // Expected: {'sum': 191, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b00011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 101,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 191, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100010; b = 8'b10011001; cin = 1'b1; // Expected: {'sum': 124, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100010; b = 8'b10011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 102,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 124, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110110; b = 8'b11000100; cin = 1'b1; // Expected: {'sum': 59, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110110; b = 8'b11000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 103,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 59, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b11001110; cin = 1'b1; // Expected: {'sum': 189, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b11001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 104,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 189, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100001; b = 8'b01001000; cin = 1'b1; // Expected: {'sum': 106, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100001; b = 8'b01001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 105,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 106, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b00100110; cin = 1'b0; // Expected: {'sum': 187, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b00100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 106,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 187, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b00010010; cin = 1'b1; // Expected: {'sum': 227, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b00010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 107,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 227, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b01110111; cin = 1'b0; // Expected: {'sum': 100, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b01110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 108,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 100, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b01010111; cin = 1'b1; // Expected: {'sum': 14, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b01010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 109,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011101; b = 8'b01011001; cin = 1'b1; // Expected: {'sum': 55, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011101; b = 8'b01011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 110,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 55, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111010; b = 8'b11100000; cin = 1'b1; // Expected: {'sum': 219, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111010; b = 8'b11100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 111,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 219, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b00100011; cin = 1'b0; // Expected: {'sum': 93, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b00100011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 112,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 93, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010111; b = 8'b11000100; cin = 1'b1; // Expected: {'sum': 28, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010111; b = 8'b11000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 113,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 28, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111011; b = 8'b01001001; cin = 1'b0; // Expected: {'sum': 196, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111011; b = 8'b01001001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 114,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 196, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b10001010; cin = 1'b0; // Expected: {'sum': 122, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b10001010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 115,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 122, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110100; b = 8'b11110111; cin = 1'b1; // Expected: {'sum': 108, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110100; b = 8'b11110111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 116,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 108, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b01111111; cin = 1'b0; // Expected: {'sum': 106, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b01111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 117,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 106, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111000; b = 8'b11101010; cin = 1'b0; // Expected: {'sum': 226, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111000; b = 8'b11101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 118,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 226, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100110; b = 8'b10101101; cin = 1'b0; // Expected: {'sum': 211, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100110; b = 8'b10101101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 119,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 211, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b10101111; cin = 1'b0; // Expected: {'sum': 240, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b10101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 120,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 240, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b01000101; cin = 1'b0; // Expected: {'sum': 212, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b01000101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 121,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 212, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111111; b = 8'b10101011; cin = 1'b1; // Expected: {'sum': 235, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111111; b = 8'b10101011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 122,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 235, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b01110010; cin = 1'b1; // Expected: {'sum': 100, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b01110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 123,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 100, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b10010100; cin = 1'b1; // Expected: {'sum': 59, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b10010100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 124,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 59, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b10100010; cin = 1'b1; // Expected: {'sum': 26, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b10100010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 125,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 26, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b00110110; cin = 1'b0; // Expected: {'sum': 63, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b00110110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 126,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 63, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b10010010; cin = 1'b1; // Expected: {'sum': 43, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b10010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 127,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 43, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b01110101; cin = 1'b0; // Expected: {'sum': 102, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b01110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 128,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 102, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b01000011; cin = 1'b0; // Expected: {'sum': 5, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b01000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 129,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 5, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b10010100; cin = 1'b0; // Expected: {'sum': 183, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b10010100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 130,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 183, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b10110000; cin = 1'b1; // Expected: {'sum': 67, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b10110000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 131,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 67, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000001; b = 8'b01010101; cin = 1'b0; // Expected: {'sum': 22, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000001; b = 8'b01010101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 132,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 22, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111001; b = 8'b10001000; cin = 1'b0; // Expected: {'sum': 193, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111001; b = 8'b10001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 133,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 193, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011110; b = 8'b11010110; cin = 1'b1; // Expected: {'sum': 181, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011110; b = 8'b11010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 134,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 181, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101000; b = 8'b01001111; cin = 1'b0; // Expected: {'sum': 119, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101000; b = 8'b01001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 135,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 119, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b11011010; cin = 1'b1; // Expected: {'sum': 253, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b11011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 136,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 253, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b11111010; cin = 1'b1; // Expected: {'sum': 14, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b11111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 137,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b00011000; cin = 1'b0; // Expected: {'sum': 74, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b00011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 138,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 74, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b10001001; cin = 1'b0; // Expected: {'sum': 135, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b10001001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 139,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 135, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b01111101; cin = 1'b0; // Expected: {'sum': 25, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b01111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 140,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 25, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001101; b = 8'b00010010; cin = 1'b1; // Expected: {'sum': 32, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001101; b = 8'b00010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 141,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 32, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b10111100; cin = 1'b1; // Expected: {'sum': 50, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b10111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 142,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 50, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010010; b = 8'b10010101; cin = 1'b1; // Expected: {'sum': 232, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010010; b = 8'b10010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 143,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 232, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b00111001; cin = 1'b0; // Expected: {'sum': 92, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b00111001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 144,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 92, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b01101111; cin = 1'b0; // Expected: {'sum': 93, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b01101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 145,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 93, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b01011101; cin = 1'b0; // Expected: {'sum': 78, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b01011101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 146,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 78, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b10110011; cin = 1'b0; // Expected: {'sum': 248, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b10110011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 147,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 248, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b00010011; cin = 1'b1; // Expected: {'sum': 152, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b00010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 148,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 152, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b00000001; cin = 1'b1; // Expected: {'sum': 147, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b00000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 149,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 147, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b00101000; cin = 1'b1; // Expected: {'sum': 209, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b00101000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 150,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 209, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b01010110; cin = 1'b0; // Expected: {'sum': 251, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b01010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 151,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 251, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100111; b = 8'b11111101; cin = 1'b1; // Expected: {'sum': 165, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100111; b = 8'b11111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 152,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 165, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b01101110; cin = 1'b0; // Expected: {'sum': 38, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b01101110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 153,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 38, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101000; b = 8'b00111010; cin = 1'b0; // Expected: {'sum': 98, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101000; b = 8'b00111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 154,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 98, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011111; b = 8'b11101111; cin = 1'b1; // Expected: {'sum': 143, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011111; b = 8'b11101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 155,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 143, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101100; b = 8'b01111111; cin = 1'b0; // Expected: {'sum': 107, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101100; b = 8'b01111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 156,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 107, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b10000101; cin = 1'b1; // Expected: {'sum': 249, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b10000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 157,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 249, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001111; b = 8'b11110011; cin = 1'b1; // Expected: {'sum': 3, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001111; b = 8'b11110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 158,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b01010110; cin = 1'b0; // Expected: {'sum': 231, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b01010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 159,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 231, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b11111001; cin = 1'b0; // Expected: {'sum': 238, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b11111001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 160,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 238, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b00111101; cin = 1'b1; // Expected: {'sum': 179, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b00111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 161,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 179, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b10100001; cin = 1'b1; // Expected: {'sum': 116, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b10100001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 162,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 116, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b00110111; cin = 1'b0; // Expected: {'sum': 109, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b00110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 163,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 109, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001100; b = 8'b01010001; cin = 1'b1; // Expected: {'sum': 30, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001100; b = 8'b01010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 164,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 30, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b11101100; cin = 1'b0; // Expected: {'sum': 117, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b11101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 165,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 117, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b11101001; cin = 1'b0; // Expected: {'sum': 215, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b11101001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 166,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 215, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b10011111; cin = 1'b1; // Expected: {'sum': 196, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b10011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 167,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 196, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101010; b = 8'b10101000; cin = 1'b1; // Expected: {'sum': 211, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101010; b = 8'b10101000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 168,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 211, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b10110100; cin = 1'b0; // Expected: {'sum': 58, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b10110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 169,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 58, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b11010011; cin = 1'b1; // Expected: {'sum': 106, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b11010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 170,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 106, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001010; b = 8'b01111101; cin = 1'b1; // Expected: {'sum': 8, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001010; b = 8'b01111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 171,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 8, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110001; b = 8'b11000110; cin = 1'b0; // Expected: {'sum': 247, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110001; b = 8'b11000110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 172,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 247, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011101; b = 8'b01010000; cin = 1'b1; // Expected: {'sum': 238, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011101; b = 8'b01010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 173,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 238, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b11110111; cin = 1'b0; // Expected: {'sum': 57, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b11110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 174,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 57, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b00001110; cin = 1'b1; // Expected: {'sum': 3, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b00001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 175,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001010; b = 8'b00100000; cin = 1'b0; // Expected: {'sum': 170, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001010; b = 8'b00100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 176,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 170, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b11011010; cin = 1'b1; // Expected: {'sum': 99, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b11011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 177,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 99, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b10101011; cin = 1'b0; // Expected: {'sum': 144, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b10101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 178,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 144, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b10000101; cin = 1'b1; // Expected: {'sum': 255, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b10000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 179,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 255, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b00110001; cin = 1'b0; // Expected: {'sum': 47, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b00110001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 180,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 47, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b01101001; cin = 1'b1; // Expected: {'sum': 160, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b01101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 181,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 160, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b01111100; cin = 1'b1; // Expected: {'sum': 20, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b01111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 182,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 20, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b11111010; cin = 1'b0; // Expected: {'sum': 207, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b11111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 183,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 207, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010111; b = 8'b00100001; cin = 1'b1; // Expected: {'sum': 121, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010111; b = 8'b00100001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 184,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 121, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b10110110; cin = 1'b1; // Expected: {'sum': 155, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b10110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 185,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 155, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001011; b = 8'b11111000; cin = 1'b1; // Expected: {'sum': 4, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001011; b = 8'b11111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 186,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010111; b = 8'b10011101; cin = 1'b1; // Expected: {'sum': 245, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010111; b = 8'b10011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 187,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 245, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b10001001; cin = 1'b1; // Expected: {'sum': 205, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b10001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 188,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 205, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100100; b = 8'b10100011; cin = 1'b0; // Expected: {'sum': 71, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100100; b = 8'b10100011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 189,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 71, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b00110010; cin = 1'b1; // Expected: {'sum': 35, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b00110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 190,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 35, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b11011001; cin = 1'b0; // Expected: {'sum': 141, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b11011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 191,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 141, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b10001010; cin = 1'b1; // Expected: {'sum': 17, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b10001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 192,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 17, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011111; b = 8'b01011010; cin = 1'b1; // Expected: {'sum': 250, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011111; b = 8'b01011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 193,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 250, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010100; b = 8'b00010111; cin = 1'b1; // Expected: {'sum': 236, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010100; b = 8'b00010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 194,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 236, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b10110000; cin = 1'b1; // Expected: {'sum': 222, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b10110000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 195,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 222, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010010; b = 8'b11111111; cin = 1'b1; // Expected: {'sum': 82, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010010; b = 8'b11111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 196,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 82, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b11010000; cin = 1'b1; // Expected: {'sum': 131, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b11010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 197,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 131, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b01110000; cin = 1'b0; // Expected: {'sum': 188, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b01110000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 198,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 188, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b10100110; cin = 1'b0; // Expected: {'sum': 188, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b10100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 199,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 188, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011111; b = 8'b01011011; cin = 1'b0; // Expected: {'sum': 250, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011111; b = 8'b01011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 200,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 250, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011010; b = 8'b10101100; cin = 1'b1; // Expected: {'sum': 7, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011010; b = 8'b10101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 201,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b11101010; cin = 1'b0; // Expected: {'sum': 28, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b11101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 202,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 28, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010001; b = 8'b00011110; cin = 1'b1; // Expected: {'sum': 240, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010001; b = 8'b00011110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 203,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 240, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b11010100; cin = 1'b0; // Expected: {'sum': 62, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b11010100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 204,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 62, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010011; b = 8'b11111111; cin = 1'b1; // Expected: {'sum': 147, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010011; b = 8'b11111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 205,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 147, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110000; b = 8'b10001001; cin = 1'b1; // Expected: {'sum': 250, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110000; b = 8'b10001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 206,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 250, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b00101000; cin = 1'b1; // Expected: {'sum': 197, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b00101000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 207,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 197, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b11101101; cin = 1'b0; // Expected: {'sum': 238, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b11101101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 208,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 238, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011100; b = 8'b10100000; cin = 1'b0; // Expected: {'sum': 124, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011100; b = 8'b10100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 209,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 124, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b01011000; cin = 1'b1; // Expected: {'sum': 65, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b01011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 210,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 65, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b10010110; cin = 1'b1; // Expected: {'sum': 38, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b10010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 211,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 38, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b10001000; cin = 1'b1; // Expected: {'sum': 118, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b10001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 212,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 118, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001010; b = 8'b01111101; cin = 1'b0; // Expected: {'sum': 7, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001010; b = 8'b01111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 213,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100010; b = 8'b00100111; cin = 1'b1; // Expected: {'sum': 10, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100010; b = 8'b00100111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 214,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b10000101; cin = 1'b1; // Expected: {'sum': 62, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b10000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 215,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 62, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110001; b = 8'b01100000; cin = 1'b1; // Expected: {'sum': 146, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110001; b = 8'b01100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 216,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 146, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001110; b = 8'b10001101; cin = 1'b0; // Expected: {'sum': 155, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001110; b = 8'b10001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 217,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 155, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101010; b = 8'b00110011; cin = 1'b1; // Expected: {'sum': 94, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101010; b = 8'b00110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 218,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 94, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101100; b = 8'b01010101; cin = 1'b1; // Expected: {'sum': 2, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101100; b = 8'b01010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 219,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b10110010; cin = 1'b1; // Expected: {'sum': 166, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b10110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 220,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 166, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010011; b = 8'b00001100; cin = 1'b0; // Expected: {'sum': 159, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010011; b = 8'b00001100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 221,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 159, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101001; b = 8'b10000111; cin = 1'b0; // Expected: {'sum': 240, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101001; b = 8'b10000111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 222,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 240, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101001; b = 8'b00001100; cin = 1'b0; // Expected: {'sum': 117, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101001; b = 8'b00001100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 223,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 117, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b01000000; cin = 1'b0; // Expected: {'sum': 93, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b01000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 224,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 93, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b10001111; cin = 1'b0; // Expected: {'sum': 124, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b10001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 225,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 124, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010101; b = 8'b00100100; cin = 1'b0; // Expected: {'sum': 57, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010101; b = 8'b00100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 226,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 57, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b01011000; cin = 1'b1; // Expected: {'sum': 17, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b01011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 227,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 17, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b00011011; cin = 1'b0; // Expected: {'sum': 27, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b00011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 228,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 27, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b01110010; cin = 1'b0; // Expected: {'sum': 24, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b01110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 229,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 24, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b11010111; cin = 1'b0; // Expected: {'sum': 89, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b11010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 230,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 89, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000101; b = 8'b01010010; cin = 1'b1; // Expected: {'sum': 24, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000101; b = 8'b01010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 231,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 24, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b00111110; cin = 1'b1; // Expected: {'sum': 104, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b00111110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 232,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 104, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101001; b = 8'b00000000; cin = 1'b1; // Expected: {'sum': 234, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101001; b = 8'b00000000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 233,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 234, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b10101111; cin = 1'b0; // Expected: {'sum': 44, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b10101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 234,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 44, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b11001110; cin = 1'b1; // Expected: {'sum': 188, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b11001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 235,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 188, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b11000111; cin = 1'b0; // Expected: {'sum': 228, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b11000111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 236,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 228, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b10011010; cin = 1'b1; // Expected: {'sum': 160, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b10011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 237,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 160, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b00110000; cin = 1'b1; // Expected: {'sum': 59, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b00110000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 238,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 59, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000111; b = 8'b11111100; cin = 1'b0; // Expected: {'sum': 131, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000111; b = 8'b11111100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 239,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 131, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b01101101; cin = 1'b0; // Expected: {'sum': 243, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b01101101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 240,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 243, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110110; b = 8'b00110100; cin = 1'b0; // Expected: {'sum': 170, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110110; b = 8'b00110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 241,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 170, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b11000111; cin = 1'b0; // Expected: {'sum': 133, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b11000111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 242,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 133, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101011; b = 8'b01001111; cin = 1'b0; // Expected: {'sum': 122, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101011; b = 8'b01001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 243,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 122, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111011; b = 8'b11001011; cin = 1'b0; // Expected: {'sum': 70, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111011; b = 8'b11001011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 244,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 70, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110011; b = 8'b11011010; cin = 1'b0; // Expected: {'sum': 141, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110011; b = 8'b11011010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 245,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 141, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111111; b = 8'b10000000; cin = 1'b1; // Expected: {'sum': 192, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111111; b = 8'b10000000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 246,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 192, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b11100011; cin = 1'b1; // Expected: {'sum': 221, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b11100011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 247,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 221, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b01011000; cin = 1'b1; // Expected: {'sum': 250, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b01011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 248,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 250, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b10101011; cin = 1'b0; // Expected: {'sum': 60, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b10101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 249,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 60, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001011; b = 8'b10011110; cin = 1'b1; // Expected: {'sum': 234, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001011; b = 8'b10011110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 250,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 234, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011011; b = 8'b10011111; cin = 1'b0; // Expected: {'sum': 186, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011011; b = 8'b10011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 251,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 186, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b10111001; cin = 1'b1; // Expected: {'sum': 49, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b10111001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 252,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 49, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b10000000; cin = 1'b0; // Expected: {'sum': 124, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b10000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 253,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 124, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b01000010; cin = 1'b1; // Expected: {'sum': 67, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b01000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 254,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 67, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010010; b = 8'b01111010; cin = 1'b1; // Expected: {'sum': 141, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010010; b = 8'b01111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 255,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 141, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b11110000; cin = 1'b1; // Expected: {'sum': 201, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b11110000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 256,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 201, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101001; b = 8'b00111101; cin = 1'b1; // Expected: {'sum': 167, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101001; b = 8'b00111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 257,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 167, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100000; b = 8'b10011001; cin = 1'b0; // Expected: {'sum': 121, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100000; b = 8'b10011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 258,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 121, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b11101001; cin = 1'b1; // Expected: {'sum': 188, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b11101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 259,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 188, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b11111100; cin = 1'b0; // Expected: {'sum': 250, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b11111100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 260,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 250, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b10010101; cin = 1'b0; // Expected: {'sum': 226, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b10010101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 261,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 226, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b11001101; cin = 1'b0; // Expected: {'sum': 64, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b11001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 262,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 64, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110110; b = 8'b10110111; cin = 1'b0; // Expected: {'sum': 45, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110110; b = 8'b10110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 263,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 45, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b10111010; cin = 1'b0; // Expected: {'sum': 179, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b10111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 264,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 179, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b10000110; cin = 1'b0; // Expected: {'sum': 234, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b10000110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 265,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 234, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011010; b = 8'b00110100; cin = 1'b1; // Expected: {'sum': 207, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011010; b = 8'b00110100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 266,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 207, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001011; b = 8'b00101010; cin = 1'b0; // Expected: {'sum': 245, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001011; b = 8'b00101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 267,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 245, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011010; b = 8'b01001001; cin = 1'b0; // Expected: {'sum': 227, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011010; b = 8'b01001001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 268,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 227, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b00101011; cin = 1'b0; // Expected: {'sum': 162, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b00101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 269,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 162, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010000; b = 8'b01100000; cin = 1'b0; // Expected: {'sum': 112, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010000; b = 8'b01100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 270,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 112, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b00010010; cin = 1'b0; // Expected: {'sum': 44, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b00010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 271,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 44, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b10110011; cin = 1'b1; // Expected: {'sum': 104, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b10110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 272,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 104, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b01011100; cin = 1'b0; // Expected: {'sum': 201, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b01011100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 273,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 201, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100110; b = 8'b11011111; cin = 1'b0; // Expected: {'sum': 197, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100110; b = 8'b11011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 274,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 197, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b01111101; cin = 1'b0; // Expected: {'sum': 44, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b01111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 275,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 44, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001110; b = 8'b11110010; cin = 1'b0; // Expected: {'sum': 64, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001110; b = 8'b11110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 276,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 64, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b11001010; cin = 1'b1; // Expected: {'sum': 233, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b11001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 277,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 233, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b00100110; cin = 1'b0; // Expected: {'sum': 198, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b00100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 278,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 198, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b01000101; cin = 1'b1; // Expected: {'sum': 241, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b01000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 279,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 241, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b10110000; cin = 1'b0; // Expected: {'sum': 122, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b10110000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 280,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 122, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000101; b = 8'b01000110; cin = 1'b0; // Expected: {'sum': 11, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000101; b = 8'b01000110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 281,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 11, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b11110000; cin = 1'b1; // Expected: {'sum': 130, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b11110000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 282,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 130, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b01111100; cin = 1'b1; // Expected: {'sum': 132, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b01111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 283,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 132, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b01001101; cin = 1'b0; // Expected: {'sum': 127, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b01001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 284,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 127, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001001; b = 8'b10000000; cin = 1'b0; // Expected: {'sum': 201, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001001; b = 8'b10000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 285,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 201, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b01111011; cin = 1'b1; // Expected: {'sum': 84, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b01111011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 286,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 84, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b10111111; cin = 1'b0; // Expected: {'sum': 28, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b10111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 287,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 28, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b00101011; cin = 1'b1; // Expected: {'sum': 63, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b00101011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 288,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 63, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100110; b = 8'b11110100; cin = 1'b0; // Expected: {'sum': 90, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100110; b = 8'b11110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 289,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 90, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001011; b = 8'b01110011; cin = 1'b0; // Expected: {'sum': 190, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001011; b = 8'b01110011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 290,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 190, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b00000111; cin = 1'b0; // Expected: {'sum': 163, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b00000111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 291,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 163, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100111; b = 8'b01101000; cin = 1'b1; // Expected: {'sum': 208, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100111; b = 8'b01101000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 292,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 208, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b11101110; cin = 1'b0; // Expected: {'sum': 166, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b11101110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 293,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 166, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b11101000; cin = 1'b1; // Expected: {'sum': 104, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b11101000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 294,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 104, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000011; b = 8'b00010011; cin = 1'b0; // Expected: {'sum': 22, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000011; b = 8'b00010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 295,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 22, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b10001001; cin = 1'b0; // Expected: {'sum': 47, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b10001001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 296,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 47, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b01100010; cin = 1'b0; // Expected: {'sum': 225, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b01100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 297,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 225, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b10011101; cin = 1'b1; // Expected: {'sum': 109, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b10011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 298,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 109, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b00101100; cin = 1'b1; // Expected: {'sum': 35, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b00101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 299,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 35, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b01011011; cin = 1'b1; // Expected: {'sum': 158, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b01011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 300,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 158, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000110; b = 8'b00011110; cin = 1'b0; // Expected: {'sum': 100, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000110; b = 8'b00011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 301,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 100, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b11111000; cin = 1'b1; // Expected: {'sum': 199, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b11111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 302,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 199, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b01110100; cin = 1'b1; // Expected: {'sum': 67, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b01110100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 303,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 67, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001011; b = 8'b01010001; cin = 1'b1; // Expected: {'sum': 93, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001011; b = 8'b01010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 304,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 93, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b01001100; cin = 1'b1; // Expected: {'sum': 108, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b01001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 305,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 108, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b11010110; cin = 1'b0; // Expected: {'sum': 138, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b11010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 306,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 138, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001101; b = 8'b00111011; cin = 1'b0; // Expected: {'sum': 8, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001101; b = 8'b00111011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 307,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 8, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b11100011; cin = 1'b1; // Expected: {'sum': 46, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b11100011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 308,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 46, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101011; b = 8'b10100110; cin = 1'b0; // Expected: {'sum': 209, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101011; b = 8'b10100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 309,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 209, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b01100111; cin = 1'b0; // Expected: {'sum': 213, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b01100111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 310,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 213, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b10011110; cin = 1'b1; // Expected: {'sum': 35, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b10011110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 311,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 35, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b01001111; cin = 1'b0; // Expected: {'sum': 223, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b01001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 312,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 223, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b00101111; cin = 1'b0; // Expected: {'sum': 186, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b00101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 313,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 186, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b00011110; cin = 1'b0; // Expected: {'sum': 249, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b00011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 314,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 249, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b10111000; cin = 1'b1; // Expected: {'sum': 53, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b10111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 315,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 53, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b11101000; cin = 1'b0; // Expected: {'sum': 41, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b11101000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 316,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 41, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b01101000; cin = 1'b0; // Expected: {'sum': 238, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b01101000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 317,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 238, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010101; b = 8'b00101001; cin = 1'b1; // Expected: {'sum': 63, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010101; b = 8'b00101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 318,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 63, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110000; b = 8'b11111011; cin = 1'b1; // Expected: {'sum': 108, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110000; b = 8'b11111011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 319,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 108, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b01100101; cin = 1'b0; // Expected: {'sum': 92, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b01100101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 320,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 92, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b10100001; cin = 1'b0; // Expected: {'sum': 24, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b10100001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 321,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 24, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011010; b = 8'b10100011; cin = 1'b1; // Expected: {'sum': 62, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011010; b = 8'b10100011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 322,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 62, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b11011111; cin = 1'b1; // Expected: {'sum': 143, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b11011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 323,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 143, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b00010011; cin = 1'b1; // Expected: {'sum': 64, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b00010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 324,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 64, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011001; b = 8'b00111101; cin = 1'b0; // Expected: {'sum': 214, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011001; b = 8'b00111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 325,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 214, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b01000111; cin = 1'b0; // Expected: {'sum': 202, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b01000111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 326,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 202, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110110; b = 8'b11001110; cin = 1'b1; // Expected: {'sum': 69, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110110; b = 8'b11001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 327,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 69, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100000; b = 8'b11011000; cin = 1'b0; // Expected: {'sum': 56, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100000; b = 8'b11011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 328,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 56, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b00100001; cin = 1'b1; // Expected: {'sum': 214, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b00100001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 329,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 214, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101100; b = 8'b01000111; cin = 1'b1; // Expected: {'sum': 52, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101100; b = 8'b01000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 330,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 52, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010100; b = 8'b01110100; cin = 1'b1; // Expected: {'sum': 201, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010100; b = 8'b01110100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 331,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 201, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110011; b = 8'b00101001; cin = 1'b0; // Expected: {'sum': 220, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110011; b = 8'b00101001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 332,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 220, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b00011110; cin = 1'b0; // Expected: {'sum': 185, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b00011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 333,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 185, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100110; b = 8'b00100001; cin = 1'b1; // Expected: {'sum': 72, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100110; b = 8'b00100001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 334,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 72, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b00111011; cin = 1'b1; // Expected: {'sum': 69, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b00111011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 335,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 69, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b01010011; cin = 1'b1; // Expected: {'sum': 20, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b01010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 336,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 20, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011010; b = 8'b10000111; cin = 1'b1; // Expected: {'sum': 34, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011010; b = 8'b10000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 337,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 34, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100110; b = 8'b01100100; cin = 1'b0; // Expected: {'sum': 74, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100110; b = 8'b01100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 338,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 74, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b01110010; cin = 1'b1; // Expected: {'sum': 75, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b01110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 339,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 75, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b11000101; cin = 1'b0; // Expected: {'sum': 77, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b11000101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 340,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 77, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b11010000; cin = 1'b0; // Expected: {'sum': 148, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b11010000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 341,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 148, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001011; b = 8'b01101001; cin = 1'b1; // Expected: {'sum': 53, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001011; b = 8'b01101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 342,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 53, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100110; b = 8'b00101010; cin = 1'b1; // Expected: {'sum': 17, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100110; b = 8'b00101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 343,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 17, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b11111110; cin = 1'b1; // Expected: {'sum': 98, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b11111110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 344,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 98, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010100; b = 8'b11111100; cin = 1'b0; // Expected: {'sum': 208, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010100; b = 8'b11111100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 345,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 208, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100010; b = 8'b01011011; cin = 1'b0; // Expected: {'sum': 253, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100010; b = 8'b01011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 346,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 253, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111000; b = 8'b10000101; cin = 1'b1; // Expected: {'sum': 190, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111000; b = 8'b10000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 347,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 190, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b11010100; cin = 1'b0; // Expected: {'sum': 106, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b11010100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 348,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 106, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b11011000; cin = 1'b1; // Expected: {'sum': 88, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b11011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 349,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 88, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011001; b = 8'b01111011; cin = 1'b1; // Expected: {'sum': 213, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011001; b = 8'b01111011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 350,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 213, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110000; b = 8'b01100010; cin = 1'b0; // Expected: {'sum': 210, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110000; b = 8'b01100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 351,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 210, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b01010110; cin = 1'b0; // Expected: {'sum': 55, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b01010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 352,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 55, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101100; b = 8'b10001000; cin = 1'b0; // Expected: {'sum': 52, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101100; b = 8'b10001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 353,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 52, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001100; b = 8'b11100000; cin = 1'b0; // Expected: {'sum': 236, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001100; b = 8'b11100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 354,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 236, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b00100101; cin = 1'b1; // Expected: {'sum': 135, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b00100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 355,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 135, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b11011000; cin = 1'b1; // Expected: {'sum': 27, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b11011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 356,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 27, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011001; b = 8'b11001101; cin = 1'b0; // Expected: {'sum': 230, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011001; b = 8'b11001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 357,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 230, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b01101010; cin = 1'b1; // Expected: {'sum': 167, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b01101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 358,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 167, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b01110110; cin = 1'b0; // Expected: {'sum': 250, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b01110110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 359,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 250, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100100; b = 8'b11101011; cin = 1'b1; // Expected: {'sum': 144, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100100; b = 8'b11101011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 360,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 144, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b00101110; cin = 1'b0; // Expected: {'sum': 183, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b00101110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 361,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 183, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110011; b = 8'b10000101; cin = 1'b1; // Expected: {'sum': 57, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110011; b = 8'b10000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 362,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 57, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b10100100; cin = 1'b1; // Expected: {'sum': 69, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b10100100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 363,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 69, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b11100100; cin = 1'b0; // Expected: {'sum': 191, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b11100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 364,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 191, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000011; b = 8'b01000111; cin = 1'b0; // Expected: {'sum': 74, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000011; b = 8'b01000111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 365,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 74, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b01000101; cin = 1'b1; // Expected: {'sum': 177, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b01000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 366,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 177, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b10001000; cin = 1'b0; // Expected: {'sum': 204, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b10001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 367,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 204, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001011; b = 8'b10000110; cin = 1'b1; // Expected: {'sum': 82, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001011; b = 8'b10000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 368,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 82, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001100; b = 8'b01110100; cin = 1'b0; // Expected: {'sum': 0, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001100; b = 8'b01110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 369,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000110; b = 8'b01100101; cin = 1'b1; // Expected: {'sum': 172, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000110; b = 8'b01100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 370,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 172, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111001; b = 8'b11000001; cin = 1'b1; // Expected: {'sum': 251, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111001; b = 8'b11000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 371,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 251, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b01001100; cin = 1'b0; // Expected: {'sum': 130, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b01001100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 372,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 130, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b10110101; cin = 1'b0; // Expected: {'sum': 217, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b10110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 373,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 217, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b10101100; cin = 1'b1; // Expected: {'sum': 159, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b10101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 374,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 159, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011010; b = 8'b00101111; cin = 1'b1; // Expected: {'sum': 10, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011010; b = 8'b00101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 375,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b10010001; cin = 1'b0; // Expected: {'sum': 147, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b10010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 376,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 147, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b00100111; cin = 1'b1; // Expected: {'sum': 138, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b00100111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 377,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 138, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b01001001; cin = 1'b0; // Expected: {'sum': 110, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b01001001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 378,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 110, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b11111011; cin = 1'b0; // Expected: {'sum': 19, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b11111011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 379,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 19, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b10000110; cin = 1'b0; // Expected: {'sum': 129, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b10000110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 380,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 129, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b00011111; cin = 1'b0; // Expected: {'sum': 3, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b00011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 381,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b01101000; cin = 1'b1; // Expected: {'sum': 92, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b01101000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 382,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 92, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b11111010; cin = 1'b1; // Expected: {'sum': 224, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b11111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 383,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 224, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b11111000; cin = 1'b1; // Expected: {'sum': 91, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b11111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 384,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 91, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b00010111; cin = 1'b0; // Expected: {'sum': 52, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b00010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 385,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 52, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b10101110; cin = 1'b1; // Expected: {'sum': 197, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b10101110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 386,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 197, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000110; b = 8'b01000101; cin = 1'b0; // Expected: {'sum': 11, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000110; b = 8'b01000101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 387,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 11, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b11110010; cin = 1'b1; // Expected: {'sum': 79, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b11110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 388,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 79, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b01111001; cin = 1'b0; // Expected: {'sum': 192, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b01111001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 389,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 192, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b11000000; cin = 1'b0; // Expected: {'sum': 36, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b11000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 390,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 36, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b10100101; cin = 1'b1; // Expected: {'sum': 147, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b10100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 391,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 147, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b01111111; cin = 1'b1; // Expected: {'sum': 18, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b01111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 392,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 18, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b11000011; cin = 1'b0; // Expected: {'sum': 94, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b11000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 393,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 94, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b00000010; cin = 1'b0; // Expected: {'sum': 25, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b00000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 394,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 25, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111000; b = 8'b00111010; cin = 1'b0; // Expected: {'sum': 50, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111000; b = 8'b00111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 395,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 50, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100000; b = 8'b01110111; cin = 1'b0; // Expected: {'sum': 87, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100000; b = 8'b01110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 396,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 87, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b01001101; cin = 1'b1; // Expected: {'sum': 186, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b01001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 397,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 186, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b11000110; cin = 1'b0; // Expected: {'sum': 18, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b11000110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 398,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 18, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b00010110; cin = 1'b1; // Expected: {'sum': 4, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b00010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 399,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b01011010; cin = 1'b1; // Expected: {'sum': 242, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b01011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 400,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 242, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000100; b = 8'b01100100; cin = 1'b0; // Expected: {'sum': 104, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000100; b = 8'b01100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 401,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 104, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b11110010; cin = 1'b1; // Expected: {'sum': 216, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b11110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 402,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 216, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b10101101; cin = 1'b0; // Expected: {'sum': 46, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b10101101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 403,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 46, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011111; b = 8'b00101110; cin = 1'b1; // Expected: {'sum': 142, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011111; b = 8'b00101110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 404,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 142, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111111; b = 8'b10111111; cin = 1'b0; // Expected: {'sum': 126, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111111; b = 8'b10111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 405,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 126, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b10001101; cin = 1'b1; // Expected: {'sum': 47, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b10001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 406,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 47, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b01100011; cin = 1'b1; // Expected: {'sum': 244, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b01100011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 407,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 244, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100010; b = 8'b10101111; cin = 1'b1; // Expected: {'sum': 146, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100010; b = 8'b10101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 408,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 146, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b00000100; cin = 1'b0; // Expected: {'sum': 9, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b00000100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 409,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 9, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b11101010; cin = 1'b0; // Expected: {'sum': 242, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b11101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 410,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 242, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b00110110; cin = 1'b1; // Expected: {'sum': 78, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b00110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 411,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 78, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b10011110; cin = 1'b1; // Expected: {'sum': 236, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b10011110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 412,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 236, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b00001001; cin = 1'b1; // Expected: {'sum': 0, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b00001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 413,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b00011101; cin = 1'b0; // Expected: {'sum': 127, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b00011101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 414,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 127, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b10101010; cin = 1'b0; // Expected: {'sum': 142, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b10101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 415,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 142, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b11111101; cin = 1'b1; // Expected: {'sum': 183, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b11111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 416,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 183, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000011; b = 8'b11111110; cin = 1'b1; // Expected: {'sum': 194, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000011; b = 8'b11111110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 417,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 194, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b00011010; cin = 1'b1; // Expected: {'sum': 93, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b00011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 418,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 93, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110000; b = 8'b10111110; cin = 1'b0; // Expected: {'sum': 46, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110000; b = 8'b10111110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 419,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 46, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110000; b = 8'b00001010; cin = 1'b1; // Expected: {'sum': 123, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110000; b = 8'b00001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 420,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 123, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b11110110; cin = 1'b1; // Expected: {'sum': 19, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b11110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 421,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 19, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001110; b = 8'b11010000; cin = 1'b0; // Expected: {'sum': 30, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001110; b = 8'b11010000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 422,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 30, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010011; b = 8'b00011000; cin = 1'b1; // Expected: {'sum': 236, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010011; b = 8'b00011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 423,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 236, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b01100111; cin = 1'b0; // Expected: {'sum': 211, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b01100111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 424,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 211, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b10111111; cin = 1'b1; // Expected: {'sum': 226, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b10111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 425,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 226, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b00101011; cin = 1'b0; // Expected: {'sum': 27, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b00101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 426,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 27, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b10001011; cin = 1'b0; // Expected: {'sum': 210, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b10001011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 427,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 210, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b01001000; cin = 1'b1; // Expected: {'sum': 193, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b01001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 428,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 193, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100010; b = 8'b01000001; cin = 1'b1; // Expected: {'sum': 36, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100010; b = 8'b01000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 429,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 36, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b00000100; cin = 1'b0; // Expected: {'sum': 206, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b00000100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 430,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 206, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b11010000; cin = 1'b0; // Expected: {'sum': 160, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b11010000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 431,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 160, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b10011001; cin = 1'b0; // Expected: {'sum': 137, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b10011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 432,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 137, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111101; b = 8'b11101101; cin = 1'b0; // Expected: {'sum': 42, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111101; b = 8'b11101101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 433,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 42, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b00001010; cin = 1'b1; // Expected: {'sum': 92, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b00001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 434,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 92, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b00011110; cin = 1'b0; // Expected: {'sum': 214, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b00011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 435,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 214, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000100; b = 8'b10101011; cin = 1'b0; // Expected: {'sum': 175, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000100; b = 8'b10101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 436,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 175, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b10001101; cin = 1'b1; // Expected: {'sum': 99, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b10001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 437,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 99, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110101; b = 8'b01000100; cin = 1'b0; // Expected: {'sum': 249, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110101; b = 8'b01000100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 438,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 249, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b11110101; cin = 1'b1; // Expected: {'sum': 7, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b11110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 439,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b11001110; cin = 1'b1; // Expected: {'sum': 100, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b11001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 440,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 100, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110011; b = 8'b11010100; cin = 1'b1; // Expected: {'sum': 136, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110011; b = 8'b11010100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 441,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 136, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100010; b = 8'b01000000; cin = 1'b0; // Expected: {'sum': 34, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100010; b = 8'b01000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 442,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 34, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b01010000; cin = 1'b0; // Expected: {'sum': 204, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b01010000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 443,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 204, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010110; b = 8'b11010000; cin = 1'b0; // Expected: {'sum': 166, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010110; b = 8'b11010000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 444,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 166, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100000; b = 8'b11011001; cin = 1'b0; // Expected: {'sum': 185, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100000; b = 8'b11011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 445,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 185, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100110; b = 8'b00101100; cin = 1'b0; // Expected: {'sum': 18, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100110; b = 8'b00101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 446,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 18, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b01001000; cin = 1'b1; // Expected: {'sum': 205, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b01001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 447,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 205, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b00000001; cin = 1'b0; // Expected: {'sum': 140, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b00000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 448,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 140, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101001; b = 8'b01010111; cin = 1'b1; // Expected: {'sum': 193, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101001; b = 8'b01010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 449,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 193, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b00100011; cin = 1'b1; // Expected: {'sum': 230, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b00100011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 450,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 230, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b10000100; cin = 1'b1; // Expected: {'sum': 174, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b10000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 451,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 174, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b10010100; cin = 1'b0; // Expected: {'sum': 108, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b10010100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 452,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 108, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b11101011; cin = 1'b0; // Expected: {'sum': 96, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b11101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 453,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 96, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001000; b = 8'b10010011; cin = 1'b1; // Expected: {'sum': 220, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001000; b = 8'b10010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 454,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 220, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001101; b = 8'b11101100; cin = 1'b0; // Expected: {'sum': 185, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001101; b = 8'b11101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 455,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 185, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b01111111; cin = 1'b0; // Expected: {'sum': 65, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b01111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 456,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 65, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101101; b = 8'b00011011; cin = 1'b1; // Expected: {'sum': 201, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101101; b = 8'b00011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 457,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 201, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111011; b = 8'b00010111; cin = 1'b0; // Expected: {'sum': 210, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111011; b = 8'b00010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 458,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 210, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b10001011; cin = 1'b0; // Expected: {'sum': 148, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b10001011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 459,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 148, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100011; b = 8'b01010110; cin = 1'b1; // Expected: {'sum': 58, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100011; b = 8'b01010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 460,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 58, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010100; b = 8'b11010001; cin = 1'b0; // Expected: {'sum': 37, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010100; b = 8'b11010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 461,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 37, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011100; b = 8'b01011110; cin = 1'b0; // Expected: {'sum': 58, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011100; b = 8'b01011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 462,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 58, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b00001101; cin = 1'b1; // Expected: {'sum': 68, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b00001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 463,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 68, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101011; b = 8'b00011000; cin = 1'b1; // Expected: {'sum': 68, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101011; b = 8'b00011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 464,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 68, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b10110110; cin = 1'b1; // Expected: {'sum': 71, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b10110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 465,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 71, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b11110000; cin = 1'b0; // Expected: {'sum': 133, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b11110000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 466,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 133, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b01001111; cin = 1'b0; // Expected: {'sum': 96, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b01001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 467,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 96, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b11011110; cin = 1'b0; // Expected: {'sum': 70, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b11011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 468,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 70, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011101; b = 8'b01011111; cin = 1'b1; // Expected: {'sum': 61, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011101; b = 8'b01011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 469,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 61, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b00111000; cin = 1'b0; // Expected: {'sum': 198, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b00111000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 470,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 198, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110011; b = 8'b00010101; cin = 1'b1; // Expected: {'sum': 201, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110011; b = 8'b00010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 471,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 201, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b00001011; cin = 1'b0; // Expected: {'sum': 196, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b00001011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 472,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 196, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b10100100; cin = 1'b1; // Expected: {'sum': 241, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b10100100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 473,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 241, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b11000001; cin = 1'b1; // Expected: {'sum': 60, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b11000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 474,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 60, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b00101111; cin = 1'b1; // Expected: {'sum': 79, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b00101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 475,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 79, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b10001000; cin = 1'b0; // Expected: {'sum': 187, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b10001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 476,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 187, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101000; b = 8'b00010001; cin = 1'b1; // Expected: {'sum': 58, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101000; b = 8'b00010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 477,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 58, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b10111110; cin = 1'b0; // Expected: {'sum': 186, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b10111110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 478,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 186, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b00000000; cin = 1'b1; // Expected: {'sum': 25, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b00000000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 479,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 25, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010011; b = 8'b11011100; cin = 1'b1; // Expected: {'sum': 112, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010011; b = 8'b11011100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 480,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 112, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b01100000; cin = 1'b0; // Expected: {'sum': 225, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b01100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 481,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 225, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111101; b = 8'b10011100; cin = 1'b0; // Expected: {'sum': 217, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111101; b = 8'b10011100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 482,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 217, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001011; b = 8'b01111111; cin = 1'b1; // Expected: {'sum': 75, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001011; b = 8'b01111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 483,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 75, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001100; b = 8'b10010010; cin = 1'b1; // Expected: {'sum': 159, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001100; b = 8'b10010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 484,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 159, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111000; b = 8'b11000000; cin = 1'b1; // Expected: {'sum': 249, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111000; b = 8'b11000000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 485,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 249, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100111; b = 8'b10110010; cin = 1'b1; // Expected: {'sum': 26, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100111; b = 8'b10110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 486,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 26, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101001; b = 8'b11000111; cin = 1'b0; // Expected: {'sum': 48, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101001; b = 8'b11000111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 487,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 48, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000011; b = 8'b00110111; cin = 1'b0; // Expected: {'sum': 58, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000011; b = 8'b00110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 488,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 58, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b01100100; cin = 1'b0; // Expected: {'sum': 204, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b01100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 489,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 204, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b01110011; cin = 1'b0; // Expected: {'sum': 100, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b01110011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 490,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 100, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b00100110; cin = 1'b1; // Expected: {'sum': 215, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b00100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 491,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 215, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b10111110; cin = 1'b1; // Expected: {'sum': 167, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b10111110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 492,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 167, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b01011100; cin = 1'b1; // Expected: {'sum': 234, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b01011100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 493,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 234, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b00010011; cin = 1'b0; // Expected: {'sum': 254, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b00010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 494,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 254, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001100; b = 8'b10010001; cin = 1'b1; // Expected: {'sum': 94, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001100; b = 8'b10010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 495,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 94, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b11101101; cin = 1'b0; // Expected: {'sum': 72, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b11101101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 496,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 72, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101111; b = 8'b00111101; cin = 1'b1; // Expected: {'sum': 45, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101111; b = 8'b00111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 497,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 45, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b10100110; cin = 1'b1; // Expected: {'sum': 86, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b10100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 498,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 86, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011010; b = 8'b00011000; cin = 1'b0; // Expected: {'sum': 242, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011010; b = 8'b00011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 499,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 242, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001001; b = 8'b01001111; cin = 1'b1; // Expected: {'sum': 25, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001001; b = 8'b01001111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 500,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 25, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b01010110; cin = 1'b1; // Expected: {'sum': 92, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b01010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 501,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 92, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010010; b = 8'b10011111; cin = 1'b1; // Expected: {'sum': 242, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010010; b = 8'b10011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 502,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 242, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101100; b = 8'b01110101; cin = 1'b0; // Expected: {'sum': 97, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101100; b = 8'b01110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 503,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 97, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b00110011; cin = 1'b1; // Expected: {'sum': 171, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b00110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 504,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 171, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b00010001; cin = 1'b1; // Expected: {'sum': 78, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b00010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 505,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 78, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b00110011; cin = 1'b1; // Expected: {'sum': 59, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b00110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 506,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 59, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b01011110; cin = 1'b0; // Expected: {'sum': 7, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b01011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 507,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011010; b = 8'b00111100; cin = 1'b0; // Expected: {'sum': 150, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011010; b = 8'b00111100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 508,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 150, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110110; b = 8'b00111100; cin = 1'b1; // Expected: {'sum': 179, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110110; b = 8'b00111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 509,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 179, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b11110101; cin = 1'b1; // Expected: {'sum': 117, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b11110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 510,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 117, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b10000110; cin = 1'b0; // Expected: {'sum': 188, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b10000110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 511,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 188, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b11011101; cin = 1'b1; // Expected: {'sum': 232, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b11011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 512,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 232, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100111; b = 8'b10111110; cin = 1'b0; // Expected: {'sum': 101, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100111; b = 8'b10111110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 513,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 101, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110001; b = 8'b00111101; cin = 1'b0; // Expected: {'sum': 174, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110001; b = 8'b00111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 514,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 174, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101110; b = 8'b00100110; cin = 1'b0; // Expected: {'sum': 84, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101110; b = 8'b00100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 515,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 84, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b01000000; cin = 1'b0; // Expected: {'sum': 186, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b01000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 516,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 186, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011010; b = 8'b11100101; cin = 1'b1; // Expected: {'sum': 64, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011010; b = 8'b11100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 517,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 64, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b11100000; cin = 1'b0; // Expected: {'sum': 37, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b11100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 518,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 37, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101111; b = 8'b10101011; cin = 1'b0; // Expected: {'sum': 218, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101111; b = 8'b10101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 519,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 218, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b01000010; cin = 1'b0; // Expected: {'sum': 116, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b01000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 520,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 116, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b01010101; cin = 1'b0; // Expected: {'sum': 206, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b01010101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 521,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 206, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b11111011; cin = 1'b1; // Expected: {'sum': 176, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b11111011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 522,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 176, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b00001010; cin = 1'b1; // Expected: {'sum': 207, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b00001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 523,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 207, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b01001000; cin = 1'b1; // Expected: {'sum': 173, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b01001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 524,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 173, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110001; b = 8'b01000001; cin = 1'b1; // Expected: {'sum': 115, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110001; b = 8'b01000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 525,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 115, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001010; b = 8'b00100100; cin = 1'b0; // Expected: {'sum': 174, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001010; b = 8'b00100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 526,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 174, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b10101011; cin = 1'b1; // Expected: {'sum': 45, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b10101011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 527,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 45, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b01010011; cin = 1'b1; // Expected: {'sum': 36, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b01010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 528,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 36, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111000; b = 8'b01001001; cin = 1'b1; // Expected: {'sum': 130, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111000; b = 8'b01001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 529,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 130, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b11111010; cin = 1'b1; // Expected: {'sum': 139, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b11111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 530,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 139, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b01011111; cin = 1'b0; // Expected: {'sum': 189, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b01011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 531,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 189, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001101; b = 8'b10011100; cin = 1'b1; // Expected: {'sum': 106, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001101; b = 8'b10011100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 532,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 106, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100000; b = 8'b00001010; cin = 1'b1; // Expected: {'sum': 43, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100000; b = 8'b00001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 533,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 43, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b01100100; cin = 1'b1; // Expected: {'sum': 198, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b01100100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 534,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 198, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b11001101; cin = 1'b0; // Expected: {'sum': 125, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b11001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 535,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 125, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110001; b = 8'b10101100; cin = 1'b1; // Expected: {'sum': 222, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110001; b = 8'b10101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 536,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 222, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b10011000; cin = 1'b0; // Expected: {'sum': 238, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b10011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 537,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 238, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b10010011; cin = 1'b1; // Expected: {'sum': 182, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b10010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 538,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 182, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b11001010; cin = 1'b1; // Expected: {'sum': 124, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b11001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 539,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 124, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b00111110; cin = 1'b1; // Expected: {'sum': 35, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b00111110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 540,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 35, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100010; b = 8'b01001010; cin = 1'b1; // Expected: {'sum': 45, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100010; b = 8'b01001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 541,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 45, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b00000011; cin = 1'b1; // Expected: {'sum': 70, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b00000011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 542,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 70, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b10100001; cin = 1'b0; // Expected: {'sum': 9, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b10100001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 543,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 9, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011010; b = 8'b01101011; cin = 1'b1; // Expected: {'sum': 70, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011010; b = 8'b01101011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 544,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 70, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b00011110; cin = 1'b1; // Expected: {'sum': 59, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b00011110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 545,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 59, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b10000010; cin = 1'b1; // Expected: {'sum': 240, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b10000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 546,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 240, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b01011101; cin = 1'b1; // Expected: {'sum': 93, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b01011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 547,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 93, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b10111000; cin = 1'b0; // Expected: {'sum': 135, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b10111000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 548,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 135, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b00010111; cin = 1'b0; // Expected: {'sum': 230, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b00010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 549,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 230, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b00111010; cin = 1'b1; // Expected: {'sum': 196, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b00111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 550,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 196, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111101; b = 8'b01110000; cin = 1'b0; // Expected: {'sum': 109, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111101; b = 8'b01110000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 551,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 109, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b10110100; cin = 1'b1; // Expected: {'sum': 107, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b10110100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 552,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 107, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b00100101; cin = 1'b1; // Expected: {'sum': 223, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b00100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 553,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 223, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b10010010; cin = 1'b0; // Expected: {'sum': 191, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b10010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 554,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 191, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100111; b = 8'b10001111; cin = 1'b0; // Expected: {'sum': 246, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100111; b = 8'b10001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 555,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 246, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000111; b = 8'b10000010; cin = 1'b1; // Expected: {'sum': 10, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000111; b = 8'b10000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 556,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111101; b = 8'b11001111; cin = 1'b1; // Expected: {'sum': 205, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111101; b = 8'b11001111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 557,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 205, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b01111000; cin = 1'b0; // Expected: {'sum': 150, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b01111000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 558,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 150, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b00000001; cin = 1'b1; // Expected: {'sum': 173, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b00000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 559,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 173, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110100; b = 8'b11101011; cin = 1'b0; // Expected: {'sum': 95, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110100; b = 8'b11101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 560,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 95, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011010; b = 8'b01001001; cin = 1'b0; // Expected: {'sum': 163, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011010; b = 8'b01001001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 561,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 163, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b00101100; cin = 1'b1; // Expected: {'sum': 253, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b00101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 562,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 253, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b00100100; cin = 1'b0; // Expected: {'sum': 21, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b00100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 563,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 21, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b11010001; cin = 1'b0; // Expected: {'sum': 218, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b11010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 564,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 218, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b01011100; cin = 1'b1; // Expected: {'sum': 157, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b01011100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 565,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 157, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010100; b = 8'b00100010; cin = 1'b0; // Expected: {'sum': 54, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010100; b = 8'b00100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 566,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 54, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b10101111; cin = 1'b1; // Expected: {'sum': 98, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b10101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 567,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 98, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111011; b = 8'b11011110; cin = 1'b1; // Expected: {'sum': 90, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111011; b = 8'b11011110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 568,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 90, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b10100101; cin = 1'b0; // Expected: {'sum': 9, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b10100101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 569,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 9, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b01111011; cin = 1'b1; // Expected: {'sum': 23, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b01111011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 570,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 23, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b11100011; cin = 1'b1; // Expected: {'sum': 3, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b11100011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 571,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b00100000; cin = 1'b0; // Expected: {'sum': 97, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b00100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 572,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 97, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b01100010; cin = 1'b0; // Expected: {'sum': 229, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b01100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 573,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 229, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b00111011; cin = 1'b1; // Expected: {'sum': 56, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b00111011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 574,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 56, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b11101000; cin = 1'b0; // Expected: {'sum': 102, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b11101000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 575,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 102, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b00101001; cin = 1'b1; // Expected: {'sum': 41, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b00101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 576,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 41, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100110; b = 8'b00001101; cin = 1'b1; // Expected: {'sum': 116, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100110; b = 8'b00001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 577,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 116, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b11100001; cin = 1'b0; // Expected: {'sum': 134, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b11100001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 578,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 134, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110001; b = 8'b00000010; cin = 1'b1; // Expected: {'sum': 52, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110001; b = 8'b00000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 579,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 52, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b00110110; cin = 1'b0; // Expected: {'sum': 239, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b00110110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 580,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 239, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000011; b = 8'b11001011; cin = 1'b0; // Expected: {'sum': 206, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000011; b = 8'b11001011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 581,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 206, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b11010000; cin = 1'b1; // Expected: {'sum': 105, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b11010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 582,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 105, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b00101011; cin = 1'b0; // Expected: {'sum': 228, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b00101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 583,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 228, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b00001110; cin = 1'b1; // Expected: {'sum': 178, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b00001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 584,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 178, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b00100110; cin = 1'b1; // Expected: {'sum': 171, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b00100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 585,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 171, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b10111001; cin = 1'b0; // Expected: {'sum': 176, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b10111001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 586,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 176, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b00010010; cin = 1'b1; // Expected: {'sum': 151, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b00010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 587,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 151, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b01011111; cin = 1'b1; // Expected: {'sum': 55, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b01011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 588,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 55, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b10110100; cin = 1'b0; // Expected: {'sum': 30, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b10110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 589,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 30, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110100; b = 8'b01001111; cin = 1'b1; // Expected: {'sum': 196, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110100; b = 8'b01001111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 590,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 196, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b00010010; cin = 1'b0; // Expected: {'sum': 14, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b00010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 591,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110111; b = 8'b00100000; cin = 1'b0; // Expected: {'sum': 87, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110111; b = 8'b00100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 592,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 87, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011111; b = 8'b01111010; cin = 1'b0; // Expected: {'sum': 217, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011111; b = 8'b01111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 593,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 217, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b01101000; cin = 1'b0; // Expected: {'sum': 94, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b01101000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 594,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 94, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001001; b = 8'b10111100; cin = 1'b1; // Expected: {'sum': 6, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001001; b = 8'b10111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 595,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101001; b = 8'b01110000; cin = 1'b1; // Expected: {'sum': 90, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101001; b = 8'b01110000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 596,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 90, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b00110100; cin = 1'b1; // Expected: {'sum': 39, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b00110100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 597,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 39, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b00110111; cin = 1'b0; // Expected: {'sum': 163, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b00110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 598,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 163, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000101; b = 8'b11001000; cin = 1'b1; // Expected: {'sum': 142, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000101; b = 8'b11001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 599,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 142, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000110; b = 8'b10010101; cin = 1'b1; // Expected: {'sum': 92, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000110; b = 8'b10010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 600,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 92, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100100; b = 8'b10100001; cin = 1'b1; // Expected: {'sum': 70, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100100; b = 8'b10100001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 601,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 70, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b10101001; cin = 1'b1; // Expected: {'sum': 244, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b10101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 602,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 244, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b10101011; cin = 1'b1; // Expected: {'sum': 74, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b10101011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 603,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 74, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b10111101; cin = 1'b1; // Expected: {'sum': 105, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b10111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 604,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 105, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111110; b = 8'b00001101; cin = 1'b0; // Expected: {'sum': 75, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111110; b = 8'b00001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 605,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 75, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b00001000; cin = 1'b0; // Expected: {'sum': 138, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b00001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 606,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 138, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b11000100; cin = 1'b1; // Expected: {'sum': 96, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b11000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 607,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 96, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000110; b = 8'b00001000; cin = 1'b1; // Expected: {'sum': 15, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000110; b = 8'b00001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 608,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101011; b = 8'b01010101; cin = 1'b0; // Expected: {'sum': 128, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101011; b = 8'b01010101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 609,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 128, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110101; b = 8'b10101111; cin = 1'b0; // Expected: {'sum': 100, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110101; b = 8'b10101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 610,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 100, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b00011001; cin = 1'b1; // Expected: {'sum': 216, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b00011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 611,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 216, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b01011010; cin = 1'b1; // Expected: {'sum': 191, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b01011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 612,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 191, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b11011000; cin = 1'b0; // Expected: {'sum': 92, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b11011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 613,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 92, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b00001110; cin = 1'b0; // Expected: {'sum': 15, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b00001110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 614,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111011; b = 8'b10011101; cin = 1'b1; // Expected: {'sum': 217, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111011; b = 8'b10011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 615,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 217, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111101; b = 8'b10000011; cin = 1'b0; // Expected: {'sum': 192, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111101; b = 8'b10000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 616,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 192, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b01110110; cin = 1'b1; // Expected: {'sum': 8, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b01110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 617,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 8, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b10111100; cin = 1'b0; // Expected: {'sum': 219, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b10111100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 618,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 219, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011101; b = 8'b11111111; cin = 1'b1; // Expected: {'sum': 157, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011101; b = 8'b11111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 619,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 157, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b00000110; cin = 1'b1; // Expected: {'sum': 43, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b00000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 620,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 43, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b10100000; cin = 1'b0; // Expected: {'sum': 196, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b10100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 621,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 196, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010111; b = 8'b11011011; cin = 1'b0; // Expected: {'sum': 50, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010111; b = 8'b11011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 622,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 50, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101101; b = 8'b10000000; cin = 1'b1; // Expected: {'sum': 46, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101101; b = 8'b10000000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 623,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 46, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000011; b = 8'b01010110; cin = 1'b1; // Expected: {'sum': 26, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000011; b = 8'b01010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 624,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 26, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000111; b = 8'b11111000; cin = 1'b1; // Expected: {'sum': 128, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000111; b = 8'b11111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 625,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 128, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b00000110; cin = 1'b1; // Expected: {'sum': 242, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b00000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 626,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 242, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b00001111; cin = 1'b1; // Expected: {'sum': 11, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b00001111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 627,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 11, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000111; b = 8'b11100100; cin = 1'b0; // Expected: {'sum': 171, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000111; b = 8'b11100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 628,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 171, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b00000100; cin = 1'b1; // Expected: {'sum': 57, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b00000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 629,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 57, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b00101010; cin = 1'b0; // Expected: {'sum': 200, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b00101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 630,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 200, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b01010010; cin = 1'b0; // Expected: {'sum': 111, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b01010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 631,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 111, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b11101111; cin = 1'b1; // Expected: {'sum': 1, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b11101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 632,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b11011100; cin = 1'b0; // Expected: {'sum': 101, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b11011100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 633,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 101, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b10001000; cin = 1'b0; // Expected: {'sum': 164, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b10001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 634,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 164, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b11100110; cin = 1'b0; // Expected: {'sum': 215, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b11100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 635,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 215, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b10111011; cin = 1'b0; // Expected: {'sum': 114, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b10111011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 636,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 114, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110000; b = 8'b11111111; cin = 1'b1; // Expected: {'sum': 112, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110000; b = 8'b11111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 637,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 112, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101010; b = 8'b01011010; cin = 1'b0; // Expected: {'sum': 132, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101010; b = 8'b01011010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 638,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 132, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b10100111; cin = 1'b1; // Expected: {'sum': 75, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b10100111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 639,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 75, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001110; b = 8'b10101000; cin = 1'b0; // Expected: {'sum': 246, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001110; b = 8'b10101000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 640,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 246, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b00111101; cin = 1'b0; // Expected: {'sum': 178, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b00111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 641,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 178, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b11101100; cin = 1'b1; // Expected: {'sum': 52, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b11101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 642,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 52, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001011; b = 8'b00100010; cin = 1'b0; // Expected: {'sum': 45, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001011; b = 8'b00100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 643,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 45, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110010; b = 8'b10111111; cin = 1'b1; // Expected: {'sum': 50, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110010; b = 8'b10111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 644,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 50, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010101; b = 8'b10010000; cin = 1'b1; // Expected: {'sum': 166, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010101; b = 8'b10010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 645,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 166, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b10100000; cin = 1'b1; // Expected: {'sum': 122, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b10100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 646,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 122, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000011; b = 8'b01100001; cin = 1'b0; // Expected: {'sum': 36, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000011; b = 8'b01100001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 647,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 36, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100110; b = 8'b01101100; cin = 1'b0; // Expected: {'sum': 82, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100110; b = 8'b01101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 648,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 82, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b10010011; cin = 1'b1; // Expected: {'sum': 254, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b10010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 649,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 254, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b00001110; cin = 1'b1; // Expected: {'sum': 197, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b00001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 650,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 197, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b00110100; cin = 1'b0; // Expected: {'sum': 51, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b00110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 651,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 51, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b00110011; cin = 1'b0; // Expected: {'sum': 243, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b00110011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 652,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 243, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b10110000; cin = 1'b1; // Expected: {'sum': 55, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b10110000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 653,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 55, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b10001100; cin = 1'b1; // Expected: {'sum': 7, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b10001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 654,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001011; b = 8'b10000001; cin = 1'b1; // Expected: {'sum': 77, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001011; b = 8'b10000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 655,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 77, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b11010100; cin = 1'b0; // Expected: {'sum': 246, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b11010100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 656,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 246, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b10001101; cin = 1'b0; // Expected: {'sum': 158, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b10001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 657,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 158, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111101; b = 8'b01010010; cin = 1'b0; // Expected: {'sum': 143, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111101; b = 8'b01010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 658,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 143, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b10110101; cin = 1'b0; // Expected: {'sum': 169, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b10110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 659,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 169, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111011; b = 8'b10111110; cin = 1'b1; // Expected: {'sum': 58, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111011; b = 8'b10111110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 660,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 58, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111111; b = 8'b11101111; cin = 1'b0; // Expected: {'sum': 46, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111111; b = 8'b11101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 661,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 46, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b10011001; cin = 1'b0; // Expected: {'sum': 41, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b10011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 662,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 41, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110111; b = 8'b10011011; cin = 1'b1; // Expected: {'sum': 211, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110111; b = 8'b10011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 663,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 211, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b00101101; cin = 1'b1; // Expected: {'sum': 44, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b00101101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 664,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 44, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b11110111; cin = 1'b0; // Expected: {'sum': 249, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b11110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 665,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 249, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110000; b = 8'b01111101; cin = 1'b1; // Expected: {'sum': 238, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110000; b = 8'b01111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 666,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 238, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b11000100; cin = 1'b0; // Expected: {'sum': 69, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b11000100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 667,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 69, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b11010110; cin = 1'b1; // Expected: {'sum': 184, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b11010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 668,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 184, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b00000001; cin = 1'b0; // Expected: {'sum': 72, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b00000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 669,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 72, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b00110001; cin = 1'b1; // Expected: {'sum': 176, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b00110001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 670,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 176, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b10101111; cin = 1'b0; // Expected: {'sum': 175, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b10101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 671,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 175, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b10001010; cin = 1'b1; // Expected: {'sum': 43, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b10001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 672,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 43, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b11001010; cin = 1'b1; // Expected: {'sum': 157, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b11001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 673,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 157, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001100; b = 8'b11010000; cin = 1'b1; // Expected: {'sum': 93, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001100; b = 8'b11010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 674,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 93, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b01001010; cin = 1'b0; // Expected: {'sum': 142, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b01001010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 675,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 142, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010100; b = 8'b10010110; cin = 1'b1; // Expected: {'sum': 43, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010100; b = 8'b10010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 676,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 43, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b00111001; cin = 1'b1; // Expected: {'sum': 218, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b00111001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 677,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 218, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010101; b = 8'b01001001; cin = 1'b1; // Expected: {'sum': 159, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010101; b = 8'b01001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 678,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 159, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b10110101; cin = 1'b0; // Expected: {'sum': 17, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b10110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 679,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 17, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000011; b = 8'b10010100; cin = 1'b1; // Expected: {'sum': 152, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000011; b = 8'b10010100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 680,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 152, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b00010010; cin = 1'b1; // Expected: {'sum': 73, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b00010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 681,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 73, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b10001000; cin = 1'b1; // Expected: {'sum': 204, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b10001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 682,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 204, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100111; b = 8'b01110111; cin = 1'b0; // Expected: {'sum': 94, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100111; b = 8'b01110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 683,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 94, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000100; b = 8'b01011001; cin = 1'b0; // Expected: {'sum': 93, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000100; b = 8'b01011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 684,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 93, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b11111010; cin = 1'b1; // Expected: {'sum': 49, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b11111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 685,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 49, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b11001010; cin = 1'b1; // Expected: {'sum': 176, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b11001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 686,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 176, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100110; b = 8'b01110010; cin = 1'b1; // Expected: {'sum': 153, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100110; b = 8'b01110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 687,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 153, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001100; b = 8'b10000001; cin = 1'b1; // Expected: {'sum': 78, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001100; b = 8'b10000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 688,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 78, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b11100100; cin = 1'b0; // Expected: {'sum': 155, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b11100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 689,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 155, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b11110100; cin = 1'b0; // Expected: {'sum': 122, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b11110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 690,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 122, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b00110101; cin = 1'b0; // Expected: {'sum': 154, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b00110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 691,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 154, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011101; b = 8'b10110000; cin = 1'b1; // Expected: {'sum': 142, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011101; b = 8'b10110000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 692,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 142, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b01011001; cin = 1'b1; // Expected: {'sum': 76, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b01011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 693,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 76, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000110; b = 8'b01011111; cin = 1'b1; // Expected: {'sum': 38, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000110; b = 8'b01011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 694,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 38, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b01001101; cin = 1'b0; // Expected: {'sum': 23, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b01001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 695,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 23, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b10110010; cin = 1'b1; // Expected: {'sum': 84, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b10110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 696,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 84, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b00010101; cin = 1'b0; // Expected: {'sum': 90, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b00010101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 697,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 90, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000101; b = 8'b10011010; cin = 1'b1; // Expected: {'sum': 96, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000101; b = 8'b10011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 698,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 96, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b10000001; cin = 1'b0; // Expected: {'sum': 113, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b10000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 699,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 113, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100111; b = 8'b10010111; cin = 1'b0; // Expected: {'sum': 190, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100111; b = 8'b10010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 700,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 190, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b01111100; cin = 1'b0; // Expected: {'sum': 5, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b01111100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 701,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 5, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100000; b = 8'b00111101; cin = 1'b0; // Expected: {'sum': 29, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100000; b = 8'b00111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 702,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 29, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b01000001; cin = 1'b0; // Expected: {'sum': 242, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b01000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 703,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 242, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b11110101; cin = 1'b1; // Expected: {'sum': 205, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b11110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 704,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 205, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b01100101; cin = 1'b0; // Expected: {'sum': 10, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b01100101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 705,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101111; b = 8'b01011011; cin = 1'b1; // Expected: {'sum': 139, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101111; b = 8'b01011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 706,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 139, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b10101000; cin = 1'b1; // Expected: {'sum': 95, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b10101000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 707,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 95, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010010; b = 8'b01011011; cin = 1'b1; // Expected: {'sum': 110, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010010; b = 8'b01011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 708,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 110, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b11000011; cin = 1'b1; // Expected: {'sum': 224, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b11000011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 709,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 224, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b00110001; cin = 1'b0; // Expected: {'sum': 40, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b00110001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 710,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 40, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b01101110; cin = 1'b1; // Expected: {'sum': 101, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b01101110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 711,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 101, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b10101101; cin = 1'b0; // Expected: {'sum': 95, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b10101101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 712,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 95, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b11111010; cin = 1'b1; // Expected: {'sum': 179, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b11111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 713,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 179, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b11101010; cin = 1'b1; // Expected: {'sum': 123, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b11101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 714,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 123, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000100; b = 8'b10111110; cin = 1'b0; // Expected: {'sum': 194, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000100; b = 8'b10111110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 715,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 194, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b11000100; cin = 1'b0; // Expected: {'sum': 66, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b11000100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 716,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 66, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b00011010; cin = 1'b1; // Expected: {'sum': 71, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b00011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 717,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 71, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b11001110; cin = 1'b1; // Expected: {'sum': 15, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b11001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 718,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010010; b = 8'b10110011; cin = 1'b0; // Expected: {'sum': 5, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010010; b = 8'b10110011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 719,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 5, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011011; b = 8'b11100010; cin = 1'b1; // Expected: {'sum': 254, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011011; b = 8'b11100010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 720,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 254, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b01111101; cin = 1'b0; // Expected: {'sum': 94, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b01111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 721,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 94, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001100; b = 8'b11101100; cin = 1'b1; // Expected: {'sum': 121, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001100; b = 8'b11101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 722,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 121, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b10000000; cin = 1'b0; // Expected: {'sum': 3, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b10000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 723,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b10101010; cin = 1'b1; // Expected: {'sum': 245, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b10101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 724,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 245, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100001; b = 8'b01000001; cin = 1'b1; // Expected: {'sum': 99, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100001; b = 8'b01000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 725,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 99, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b11111111; cin = 1'b0; // Expected: {'sum': 209, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b11111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 726,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 209, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101110; b = 8'b01010010; cin = 1'b1; // Expected: {'sum': 1, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101110; b = 8'b01010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 727,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b00111000; cin = 1'b0; // Expected: {'sum': 2, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b00111000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 728,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011011; b = 8'b10011100; cin = 1'b0; // Expected: {'sum': 183, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011011; b = 8'b10011100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 729,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 183, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000111; b = 8'b10001110; cin = 1'b1; // Expected: {'sum': 22, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000111; b = 8'b10001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 730,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 22, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010100; b = 8'b01101111; cin = 1'b1; // Expected: {'sum': 196, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010100; b = 8'b01101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 731,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 196, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b11001011; cin = 1'b0; // Expected: {'sum': 28, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b11001011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 732,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 28, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b11100010; cin = 1'b0; // Expected: {'sum': 119, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b11100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 733,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 119, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b01100000; cin = 1'b1; // Expected: {'sum': 252, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b01100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 734,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 252, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b01011010; cin = 1'b0; // Expected: {'sum': 113, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b01011010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 735,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 113, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b11110110; cin = 1'b0; // Expected: {'sum': 34, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b11110110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 736,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 34, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b10010010; cin = 1'b0; // Expected: {'sum': 255, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b10010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 737,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 255, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111111; b = 8'b01010000; cin = 1'b1; // Expected: {'sum': 144, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111111; b = 8'b01010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 738,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 144, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b00001100; cin = 1'b1; // Expected: {'sum': 184, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b00001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 739,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 184, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101101; b = 8'b00101010; cin = 1'b0; // Expected: {'sum': 215, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101101; b = 8'b00101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 740,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 215, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100111; b = 8'b01010001; cin = 1'b0; // Expected: {'sum': 120, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100111; b = 8'b01010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 741,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 120, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b10001001; cin = 1'b0; // Expected: {'sum': 88, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b10001001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 742,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 88, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b01001011; cin = 1'b0; // Expected: {'sum': 225, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b01001011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 743,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 225, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001111; b = 8'b11000010; cin = 1'b0; // Expected: {'sum': 209, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001111; b = 8'b11000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 744,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 209, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b10011111; cin = 1'b0; // Expected: {'sum': 27, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b10011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 745,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 27, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110000; b = 8'b01110111; cin = 1'b1; // Expected: {'sum': 232, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110000; b = 8'b01110111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 746,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 232, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b00010100; cin = 1'b1; // Expected: {'sum': 98, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b00010100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 747,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 98, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b11010100; cin = 1'b0; // Expected: {'sum': 234, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b11010100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 748,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 234, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b10111111; cin = 1'b0; // Expected: {'sum': 215, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b10111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 749,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 215, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110011; b = 8'b11000101; cin = 1'b1; // Expected: {'sum': 121, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110011; b = 8'b11000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 750,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 121, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b01101010; cin = 1'b1; // Expected: {'sum': 188, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b01101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 751,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 188, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b01110100; cin = 1'b0; // Expected: {'sum': 231, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b01110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 752,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 231, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b01011010; cin = 1'b0; // Expected: {'sum': 74, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b01011010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 753,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 74, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101010; b = 8'b11011110; cin = 1'b0; // Expected: {'sum': 8, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101010; b = 8'b11011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 754,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 8, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b00100111; cin = 1'b0; // Expected: {'sum': 143, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b00100111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 755,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 143, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010000; b = 8'b10010111; cin = 1'b1; // Expected: {'sum': 168, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010000; b = 8'b10010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 756,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 168, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b11001100; cin = 1'b1; // Expected: {'sum': 90, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b11001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 757,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 90, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b00001001; cin = 1'b1; // Expected: {'sum': 64, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b00001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 758,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 64, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010111; b = 8'b11101100; cin = 1'b0; // Expected: {'sum': 67, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010111; b = 8'b11101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 759,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 67, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b11001101; cin = 1'b0; // Expected: {'sum': 177, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b11001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 760,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 177, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b01010011; cin = 1'b1; // Expected: {'sum': 18, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b01010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 761,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 18, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b01100001; cin = 1'b0; // Expected: {'sum': 85, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b01100001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 762,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 85, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b10001011; cin = 1'b1; // Expected: {'sum': 103, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b10001011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 763,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 103, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001101; b = 8'b01111111; cin = 1'b0; // Expected: {'sum': 140, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001101; b = 8'b01111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 764,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 140, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111011; b = 8'b11111001; cin = 1'b1; // Expected: {'sum': 53, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111011; b = 8'b11111001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 765,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 53, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b01110110; cin = 1'b1; // Expected: {'sum': 46, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b01110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 766,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 46, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100001; b = 8'b10011001; cin = 1'b1; // Expected: {'sum': 187, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100001; b = 8'b10011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 767,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 187, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b11000010; cin = 1'b0; // Expected: {'sum': 248, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b11000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 768,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 248, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011010; b = 8'b01010001; cin = 1'b0; // Expected: {'sum': 171, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011010; b = 8'b01010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 769,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 171, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010001; b = 8'b10010100; cin = 1'b1; // Expected: {'sum': 102, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010001; b = 8'b10010100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 770,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 102, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b11011010; cin = 1'b0; // Expected: {'sum': 131, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b11011010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 771,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 131, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b00110001; cin = 1'b0; // Expected: {'sum': 68, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b00110001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 772,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 68, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b10011100; cin = 1'b1; // Expected: {'sum': 249, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b10011100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 773,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 249, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b01011011; cin = 1'b0; // Expected: {'sum': 199, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b01011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 774,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 199, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b11100011; cin = 1'b1; // Expected: {'sum': 201, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b11100011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 775,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 201, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b11000001; cin = 1'b1; // Expected: {'sum': 96, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b11000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 776,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 96, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b10110010; cin = 1'b0; // Expected: {'sum': 246, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b10110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 777,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 246, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011101; b = 8'b00000010; cin = 1'b1; // Expected: {'sum': 224, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011101; b = 8'b00000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 778,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 224, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b00111100; cin = 1'b0; // Expected: {'sum': 243, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b00111100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 779,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 243, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b00010010; cin = 1'b0; // Expected: {'sum': 119, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b00010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 780,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 119, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110110; b = 8'b01111111; cin = 1'b0; // Expected: {'sum': 245, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110110; b = 8'b01111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 781,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 245, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b00111011; cin = 1'b0; // Expected: {'sum': 38, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b00111011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 782,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 38, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100010; b = 8'b01000001; cin = 1'b0; // Expected: {'sum': 35, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100010; b = 8'b01000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 783,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 35, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010011; b = 8'b00110100; cin = 1'b1; // Expected: {'sum': 136, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010011; b = 8'b00110100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 784,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 136, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111111; b = 8'b11100000; cin = 1'b1; // Expected: {'sum': 160, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111111; b = 8'b11100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 785,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 160, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b10010000; cin = 1'b1; // Expected: {'sum': 74, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b10010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 786,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 74, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b10000111; cin = 1'b0; // Expected: {'sum': 244, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b10000111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 787,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 244, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b01101110; cin = 1'b0; // Expected: {'sum': 227, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b01101110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 788,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 227, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b01011111; cin = 1'b1; // Expected: {'sum': 87, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b01011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 789,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 87, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011001; b = 8'b10011001; cin = 1'b0; // Expected: {'sum': 50, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011001; b = 8'b10011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 790,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 50, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b00100000; cin = 1'b0; // Expected: {'sum': 139, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b00100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 791,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 139, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b10001110; cin = 1'b1; // Expected: {'sum': 81, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b10001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 792,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 81, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b10111001; cin = 1'b0; // Expected: {'sum': 174, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b10111001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 793,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 174, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b11110011; cin = 1'b1; // Expected: {'sum': 24, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b11110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 794,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 24, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b00111000; cin = 1'b0; // Expected: {'sum': 177, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b00111000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 795,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 177, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b11010000; cin = 1'b1; // Expected: {'sum': 60, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b11010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 796,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 60, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101100; b = 8'b01111100; cin = 1'b0; // Expected: {'sum': 40, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101100; b = 8'b01111100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 797,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 40, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011111; b = 8'b00000100; cin = 1'b1; // Expected: {'sum': 100, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011111; b = 8'b00000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 798,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 100, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010000; b = 8'b01000101; cin = 1'b1; // Expected: {'sum': 86, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010000; b = 8'b01000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 799,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 86, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b11000001; cin = 1'b0; // Expected: {'sum': 52, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b11000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 800,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 52, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b10001000; cin = 1'b1; // Expected: {'sum': 159, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b10001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 801,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 159, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b10000011; cin = 1'b0; // Expected: {'sum': 197, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b10000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 802,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 197, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b11010001; cin = 1'b1; // Expected: {'sum': 244, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b11010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 803,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 244, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b10111111; cin = 1'b0; // Expected: {'sum': 0, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b10111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 804,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111110; b = 8'b10001111; cin = 1'b1; // Expected: {'sum': 206, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111110; b = 8'b10001111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 805,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 206, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b01111010; cin = 1'b1; // Expected: {'sum': 107, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b01111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 806,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 107, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b11010111; cin = 1'b1; // Expected: {'sum': 188, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b11010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 807,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 188, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b01100001; cin = 1'b1; // Expected: {'sum': 128, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b01100001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 808,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 128, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b01011010; cin = 1'b1; // Expected: {'sum': 235, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b01011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 809,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 235, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b11011001; cin = 1'b1; // Expected: {'sum': 142, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b11011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 810,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 142, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011111; b = 8'b00100110; cin = 1'b0; // Expected: {'sum': 197, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011111; b = 8'b00100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 811,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 197, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001100; b = 8'b00010000; cin = 1'b1; // Expected: {'sum': 221, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001100; b = 8'b00010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 812,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 221, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b10011010; cin = 1'b0; // Expected: {'sum': 111, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b10011010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 813,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 111, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110000; b = 8'b01110000; cin = 1'b1; // Expected: {'sum': 161, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110000; b = 8'b01110000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 814,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 161, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b10101100; cin = 1'b1; // Expected: {'sum': 202, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b10101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 815,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 202, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110000; b = 8'b01011000; cin = 1'b1; // Expected: {'sum': 201, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110000; b = 8'b01011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 816,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 201, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100100; b = 8'b11110110; cin = 1'b0; // Expected: {'sum': 154, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100100; b = 8'b11110110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 817,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 154, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b11101000; cin = 1'b0; // Expected: {'sum': 208, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b11101000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 818,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 208, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b11000000; cin = 1'b1; // Expected: {'sum': 172, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b11000000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 819,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 172, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b11010011; cin = 1'b0; // Expected: {'sum': 161, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b11010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 820,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 161, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b01101100; cin = 1'b1; // Expected: {'sum': 30, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b01101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 821,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 30, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111011; b = 8'b10001010; cin = 1'b1; // Expected: {'sum': 198, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111011; b = 8'b10001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 822,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 198, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b10011111; cin = 1'b0; // Expected: {'sum': 240, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b10011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 823,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 240, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b01001110; cin = 1'b1; // Expected: {'sum': 179, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b01001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 824,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 179, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b00000011; cin = 1'b0; // Expected: {'sum': 94, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b00000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 825,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 94, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101001; b = 8'b00001110; cin = 1'b1; // Expected: {'sum': 120, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101001; b = 8'b00001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 826,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 120, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b00111010; cin = 1'b0; // Expected: {'sum': 51, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b00111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 827,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 51, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b01111010; cin = 1'b1; // Expected: {'sum': 86, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b01111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 828,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 86, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b01101111; cin = 1'b1; // Expected: {'sum': 244, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b01101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 829,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 244, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b01011111; cin = 1'b0; // Expected: {'sum': 203, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b01011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 830,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 203, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b10110101; cin = 1'b0; // Expected: {'sum': 19, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b10110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 831,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 19, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b01100000; cin = 1'b0; // Expected: {'sum': 220, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b01100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 832,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 220, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001101; b = 8'b00101100; cin = 1'b1; // Expected: {'sum': 58, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001101; b = 8'b00101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 833,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 58, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101010; b = 8'b01011110; cin = 1'b0; // Expected: {'sum': 8, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101010; b = 8'b01011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 834,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 8, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100111; b = 8'b01000110; cin = 1'b1; // Expected: {'sum': 46, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100111; b = 8'b01000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 835,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 46, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101011; b = 8'b01101101; cin = 1'b0; // Expected: {'sum': 152, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101011; b = 8'b01101101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 836,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 152, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000111; b = 8'b11000001; cin = 1'b1; // Expected: {'sum': 137, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000111; b = 8'b11000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 837,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 137, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b01001101; cin = 1'b0; // Expected: {'sum': 87, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b01001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 838,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 87, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b11111100; cin = 1'b0; // Expected: {'sum': 4, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b11111100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 839,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b11001001; cin = 1'b1; // Expected: {'sum': 228, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b11001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 840,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 228, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110001; b = 8'b01000100; cin = 1'b1; // Expected: {'sum': 118, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110001; b = 8'b01000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 841,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 118, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110110; b = 8'b11100110; cin = 1'b0; // Expected: {'sum': 92, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110110; b = 8'b11100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 842,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 92, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b01010001; cin = 1'b1; // Expected: {'sum': 22, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b01010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 843,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 22, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b11110011; cin = 1'b1; // Expected: {'sum': 115, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b11110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 844,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 115, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b01111111; cin = 1'b1; // Expected: {'sum': 33, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b01111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 845,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 33, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b01100011; cin = 1'b1; // Expected: {'sum': 76, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b01100011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 846,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 76, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110000; b = 8'b01110000; cin = 1'b0; // Expected: {'sum': 160, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110000; b = 8'b01110000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 847,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 160, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010100; b = 8'b01110100; cin = 1'b0; // Expected: {'sum': 8, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010100; b = 8'b01110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 848,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 8, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b01000001; cin = 1'b0; // Expected: {'sum': 146, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b01000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 849,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 146, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000101; b = 8'b10000011; cin = 1'b1; // Expected: {'sum': 9, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000101; b = 8'b10000011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 850,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 9, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010011; b = 8'b01010011; cin = 1'b1; // Expected: {'sum': 231, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010011; b = 8'b01010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 851,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 231, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010101; b = 8'b10111100; cin = 1'b0; // Expected: {'sum': 209, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010101; b = 8'b10111100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 852,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 209, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b00110101; cin = 1'b1; // Expected: {'sum': 76, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b00110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 853,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 76, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b00010101; cin = 1'b0; // Expected: {'sum': 145, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b00010101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 854,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 145, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b00111101; cin = 1'b1; // Expected: {'sum': 52, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b00111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 855,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 52, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b01111000; cin = 1'b1; // Expected: {'sum': 166, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b01111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 856,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 166, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b01010110; cin = 1'b0; // Expected: {'sum': 75, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b01010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 857,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 75, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b10011110; cin = 1'b0; // Expected: {'sum': 249, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b10011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 858,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 249, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b00111011; cin = 1'b0; // Expected: {'sum': 201, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b00111011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 859,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 201, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b11100001; cin = 1'b0; // Expected: {'sum': 13, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b11100001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 860,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 13, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b11000100; cin = 1'b0; // Expected: {'sum': 224, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b11000100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 861,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 224, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001001; b = 8'b01011000; cin = 1'b1; // Expected: {'sum': 34, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001001; b = 8'b01011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 862,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 34, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b11111111; cin = 1'b0; // Expected: {'sum': 103, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b11111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 863,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 103, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b10000100; cin = 1'b1; // Expected: {'sum': 241, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b10000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 864,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 241, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b00111011; cin = 1'b1; // Expected: {'sum': 189, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b00111011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 865,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 189, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b10101111; cin = 1'b0; // Expected: {'sum': 29, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b10101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 866,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 29, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001011; b = 8'b01101010; cin = 1'b1; // Expected: {'sum': 118, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001011; b = 8'b01101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 867,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 118, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b11010001; cin = 1'b1; // Expected: {'sum': 169, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b11010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 868,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 169, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b00110010; cin = 1'b1; // Expected: {'sum': 237, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b00110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 869,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 237, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b01010110; cin = 1'b0; // Expected: {'sum': 59, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b01010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 870,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 59, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b01101100; cin = 1'b0; // Expected: {'sum': 80, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b01101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 871,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 80, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b01111011; cin = 1'b1; // Expected: {'sum': 243, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b01111011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 872,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 243, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b00001101; cin = 1'b1; // Expected: {'sum': 58, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b00001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 873,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 58, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b01110001; cin = 1'b1; // Expected: {'sum': 246, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b01110001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 874,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 246, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110010; b = 8'b00011111; cin = 1'b1; // Expected: {'sum': 146, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110010; b = 8'b00011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 875,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 146, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b10011110; cin = 1'b0; // Expected: {'sum': 166, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b10011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 876,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 166, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111111; b = 8'b01000110; cin = 1'b0; // Expected: {'sum': 5, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111111; b = 8'b01000110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 877,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 5, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b01010000; cin = 1'b0; // Expected: {'sum': 102, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b01010000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 878,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 102, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b00011110; cin = 1'b0; // Expected: {'sum': 155, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b00011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 879,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 155, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100111; b = 8'b10111011; cin = 1'b0; // Expected: {'sum': 226, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100111; b = 8'b10111011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 880,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 226, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b11110100; cin = 1'b0; // Expected: {'sum': 22, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b11110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 881,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 22, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b10100100; cin = 1'b1; // Expected: {'sum': 15, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b10100100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 882,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b00110001; cin = 1'b0; // Expected: {'sum': 231, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b00110001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 883,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 231, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b11011111; cin = 1'b0; // Expected: {'sum': 224, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b11011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 884,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 224, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100111; b = 8'b00011011; cin = 1'b1; // Expected: {'sum': 131, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100111; b = 8'b00011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 885,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 131, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b10110000; cin = 1'b0; // Expected: {'sum': 135, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b10110000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 886,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 135, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b01001011; cin = 1'b1; // Expected: {'sum': 252, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b01001011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 887,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 252, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b00111110; cin = 1'b0; // Expected: {'sum': 192, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b00111110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 888,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 192, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b11110010; cin = 1'b1; // Expected: {'sum': 248, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b11110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 889,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 248, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111101; b = 8'b00101100; cin = 1'b0; // Expected: {'sum': 105, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111101; b = 8'b00101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 890,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 105, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000100; b = 8'b00000111; cin = 1'b1; // Expected: {'sum': 12, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000100; b = 8'b00000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 891,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 12, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011001; b = 8'b10011000; cin = 1'b0; // Expected: {'sum': 49, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011001; b = 8'b10011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 892,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 49, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101001; b = 8'b00101111; cin = 1'b0; // Expected: {'sum': 152, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101001; b = 8'b00101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 893,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 152, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b00011011; cin = 1'b0; // Expected: {'sum': 85, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b00011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 894,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 85, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010001; b = 8'b10100001; cin = 1'b0; // Expected: {'sum': 114, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010001; b = 8'b10100001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 895,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 114, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b01110010; cin = 1'b1; // Expected: {'sum': 245, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b01110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 896,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 245, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111110; b = 8'b00000010; cin = 1'b1; // Expected: {'sum': 65, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111110; b = 8'b00000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 897,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 65, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b10000010; cin = 1'b0; // Expected: {'sum': 68, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b10000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 898,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 68, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b11011110; cin = 1'b0; // Expected: {'sum': 87, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b11011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 899,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 87, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100010; b = 8'b00101011; cin = 1'b0; // Expected: {'sum': 13, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100010; b = 8'b00101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 900,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 13, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b10011000; cin = 1'b1; // Expected: {'sum': 34, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b10011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 901,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 34, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011101; b = 8'b01110011; cin = 1'b1; // Expected: {'sum': 81, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011101; b = 8'b01110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 902,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 81, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011101; b = 8'b01011010; cin = 1'b1; // Expected: {'sum': 56, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011101; b = 8'b01011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 903,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 56, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b10101010; cin = 1'b0; // Expected: {'sum': 106, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b10101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 904,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 106, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b11110111; cin = 1'b0; // Expected: {'sum': 84, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b11110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 905,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 84, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b11001101; cin = 1'b1; // Expected: {'sum': 99, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b11001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 906,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 99, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100111; b = 8'b11110000; cin = 1'b1; // Expected: {'sum': 24, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100111; b = 8'b11110000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 907,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 24, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111101; b = 8'b10110110; cin = 1'b0; // Expected: {'sum': 243, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111101; b = 8'b10110110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 908,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 243, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b10000100; cin = 1'b1; // Expected: {'sum': 9, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b10000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 909,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 9, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b01000110; cin = 1'b1; // Expected: {'sum': 197, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b01000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 910,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 197, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001101; b = 8'b11101100; cin = 1'b1; // Expected: {'sum': 250, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001101; b = 8'b11101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 911,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 250, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b10000001; cin = 1'b1; // Expected: {'sum': 59, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b10000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 912,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 59, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111101; b = 8'b01101011; cin = 1'b1; // Expected: {'sum': 169, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111101; b = 8'b01101011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 913,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 169, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b11100001; cin = 1'b0; // Expected: {'sum': 10, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b11100001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 914,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b10000111; cin = 1'b0; // Expected: {'sum': 108, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b10000111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 915,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 108, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b11100010; cin = 1'b0; // Expected: {'sum': 158, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b11100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 916,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 158, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011111; b = 8'b11001110; cin = 1'b1; // Expected: {'sum': 46, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011111; b = 8'b11001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 917,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 46, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b00000100; cin = 1'b0; // Expected: {'sum': 196, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b00000100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 918,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 196, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101001; b = 8'b11100010; cin = 1'b1; // Expected: {'sum': 204, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101001; b = 8'b11100010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 919,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 204, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b11000101; cin = 1'b0; // Expected: {'sum': 173, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b11000101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 920,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 173, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b00101101; cin = 1'b1; // Expected: {'sum': 55, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b00101101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 921,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 55, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b11010001; cin = 1'b1; // Expected: {'sum': 198, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b11010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 922,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 198, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100011; b = 8'b11110010; cin = 1'b0; // Expected: {'sum': 213, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100011; b = 8'b11110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 923,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 213, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b00011101; cin = 1'b0; // Expected: {'sum': 109, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b00011101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 924,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 109, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000111; b = 8'b10110010; cin = 1'b0; // Expected: {'sum': 121, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000111; b = 8'b10110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 925,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 121, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b11110111; cin = 1'b0; // Expected: {'sum': 242, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b11110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 926,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 242, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b10101110; cin = 1'b0; // Expected: {'sum': 76, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b10101110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 927,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 76, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b00111011; cin = 1'b0; // Expected: {'sum': 159, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b00111011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 928,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 159, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b11000110; cin = 1'b0; // Expected: {'sum': 206, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b11000110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 929,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 206, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b10001101; cin = 1'b1; // Expected: {'sum': 124, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b10001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 930,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 124, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b01111010; cin = 1'b0; // Expected: {'sum': 237, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b01111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 931,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 237, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b00000001; cin = 1'b0; // Expected: {'sum': 53, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b00000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 932,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 53, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b10011010; cin = 1'b0; // Expected: {'sum': 245, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b10011010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 933,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 245, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b01001001; cin = 1'b0; // Expected: {'sum': 54, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b01001001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 934,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 54, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b00010011; cin = 1'b0; // Expected: {'sum': 17, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b00010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 935,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 17, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b00101010; cin = 1'b1; // Expected: {'sum': 187, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b00101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 936,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 187, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110001; b = 8'b11000100; cin = 1'b0; // Expected: {'sum': 53, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110001; b = 8'b11000100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 937,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 53, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b10110111; cin = 1'b1; // Expected: {'sum': 21, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b10110111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 938,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 21, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b00110100; cin = 1'b1; // Expected: {'sum': 127, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b00110100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 939,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 127, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b10110001; cin = 1'b0; // Expected: {'sum': 1, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b10110001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 940,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011100; b = 8'b10001000; cin = 1'b1; // Expected: {'sum': 101, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011100; b = 8'b10001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 941,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 101, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b10111001; cin = 1'b0; // Expected: {'sum': 146, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b10111001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 942,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 146, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110001; b = 8'b11111100; cin = 1'b0; // Expected: {'sum': 109, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110001; b = 8'b11111100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 943,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 109, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b10111101; cin = 1'b1; // Expected: {'sum': 142, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b10111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 944,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 142, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b01000100; cin = 1'b0; // Expected: {'sum': 175, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b01000100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 945,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 175, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010101; b = 8'b10110110; cin = 1'b1; // Expected: {'sum': 12, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010101; b = 8'b10110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 946,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010100; b = 8'b01111011; cin = 1'b0; // Expected: {'sum': 207, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010100; b = 8'b01111011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 947,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 207, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b01011101; cin = 1'b1; // Expected: {'sum': 46, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b01011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 948,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 46, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101110; b = 8'b10100111; cin = 1'b0; // Expected: {'sum': 85, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101110; b = 8'b10100111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 949,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 85, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b11010011; cin = 1'b1; // Expected: {'sum': 85, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b11010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 950,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 85, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b11100101; cin = 1'b1; // Expected: {'sum': 180, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b11100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 951,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 180, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110010; b = 8'b00101110; cin = 1'b0; // Expected: {'sum': 160, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110010; b = 8'b00101110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 952,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 160, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101001; b = 8'b10100110; cin = 1'b0; // Expected: {'sum': 15, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101001; b = 8'b10100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 953,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b10111111; cin = 1'b1; // Expected: {'sum': 68, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b10111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 954,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 68, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b01001011; cin = 1'b1; // Expected: {'sum': 2, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b01001011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 955,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111001; b = 8'b10101100; cin = 1'b1; // Expected: {'sum': 230, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111001; b = 8'b10101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 956,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 230, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b00001101; cin = 1'b1; // Expected: {'sum': 42, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b00001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 957,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 42, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b10001010; cin = 1'b0; // Expected: {'sum': 42, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b10001010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 958,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 42, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101100; b = 8'b10001011; cin = 1'b0; // Expected: {'sum': 119, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101100; b = 8'b10001011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 959,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 119, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b11010100; cin = 1'b0; // Expected: {'sum': 66, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b11010100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 960,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 66, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b11001110; cin = 1'b0; // Expected: {'sum': 14, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b11001110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 961,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001101; b = 8'b11100110; cin = 1'b1; // Expected: {'sum': 244, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001101; b = 8'b11100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 962,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 244, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000011; b = 8'b01011011; cin = 1'b1; // Expected: {'sum': 31, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000011; b = 8'b01011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 963,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 31, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b00000001; cin = 1'b0; // Expected: {'sum': 246, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b00000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 964,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 246, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b10111101; cin = 1'b1; // Expected: {'sum': 3, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b10111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 965,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001101; b = 8'b10101011; cin = 1'b0; // Expected: {'sum': 184, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001101; b = 8'b10101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 966,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 184, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b00000011; cin = 1'b0; // Expected: {'sum': 4, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b00000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 967,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 4, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b00001011; cin = 1'b0; // Expected: {'sum': 69, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b00001011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 968,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 69, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b00110011; cin = 1'b1; // Expected: {'sum': 169, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b00110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 969,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 169, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b00000011; cin = 1'b0; // Expected: {'sum': 37, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b00000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 970,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 37, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b11101010; cin = 1'b0; // Expected: {'sum': 180, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b11101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 971,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 180, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010011; b = 8'b01011011; cin = 1'b1; // Expected: {'sum': 175, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010011; b = 8'b01011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 972,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 175, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111011; b = 8'b01011100; cin = 1'b0; // Expected: {'sum': 23, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111011; b = 8'b01011100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 973,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 23, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b10110111; cin = 1'b1; // Expected: {'sum': 32, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b10110111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 974,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 32, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b00110110; cin = 1'b1; // Expected: {'sum': 106, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b00110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 975,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 106, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001101; b = 8'b01111110; cin = 1'b0; // Expected: {'sum': 75, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001101; b = 8'b01111110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 976,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 75, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b01000100; cin = 1'b0; // Expected: {'sum': 109, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b01000100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 977,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 109, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b10011111; cin = 1'b0; // Expected: {'sum': 87, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b10011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 978,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 87, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b10101011; cin = 1'b0; // Expected: {'sum': 159, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b10101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 979,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 159, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101000; b = 8'b10110010; cin = 1'b1; // Expected: {'sum': 219, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101000; b = 8'b10110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 980,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 219, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b10000011; cin = 1'b0; // Expected: {'sum': 162, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b10000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 981,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 162, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101110; b = 8'b11100000; cin = 1'b0; // Expected: {'sum': 14, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101110; b = 8'b11100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 982,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b01110010; cin = 1'b0; // Expected: {'sum': 188, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b01110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 983,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 188, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b00011010; cin = 1'b0; // Expected: {'sum': 124, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b00011010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 984,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 124, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b00000111; cin = 1'b1; // Expected: {'sum': 76, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b00000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 985,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 76, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011111; b = 8'b10000000; cin = 1'b1; // Expected: {'sum': 32, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011111; b = 8'b10000000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 986,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 32, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110000; b = 8'b00000110; cin = 1'b1; // Expected: {'sum': 119, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110000; b = 8'b00000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 987,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 119, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b01001000; cin = 1'b0; // Expected: {'sum': 33, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b01001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 988,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 33, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b01111000; cin = 1'b0; // Expected: {'sum': 30, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b01111000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 989,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 30, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b00111110; cin = 1'b0; // Expected: {'sum': 177, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b00111110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 990,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 177, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100110; b = 8'b01000101; cin = 1'b1; // Expected: {'sum': 108, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100110; b = 8'b01000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 991,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 108, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b11100111; cin = 1'b0; // Expected: {'sum': 20, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b11100111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 992,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 20, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001011; b = 8'b01010000; cin = 1'b1; // Expected: {'sum': 92, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001011; b = 8'b01010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 993,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 92, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b00000101; cin = 1'b0; // Expected: {'sum': 242, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b00000101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 994,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 242, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111011; b = 8'b00100010; cin = 1'b0; // Expected: {'sum': 157, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111011; b = 8'b00100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 995,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 157, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b00011010; cin = 1'b0; // Expected: {'sum': 189, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b00011010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 996,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 189, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b01110101; cin = 1'b0; // Expected: {'sum': 253, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b01110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 997,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 253, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b11010100; cin = 1'b0; // Expected: {'sum': 220, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b11010100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 998,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 220, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111111; b = 8'b10011001; cin = 1'b1; // Expected: {'sum': 217, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111111; b = 8'b10011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 999,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 217, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001000; b = 8'b10000011; cin = 1'b0; // Expected: {'sum': 203, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001000; b = 8'b10000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1000,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 203, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b01101111; cin = 1'b1; // Expected: {'sum': 189, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b01101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1001,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 189, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100010; b = 8'b11111001; cin = 1'b1; // Expected: {'sum': 156, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100010; b = 8'b11111001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1002,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 156, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b11000110; cin = 1'b0; // Expected: {'sum': 33, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b11000110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1003,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 33, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b10000000; cin = 1'b1; // Expected: {'sum': 62, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b10000000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1004,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 62, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b01011000; cin = 1'b0; // Expected: {'sum': 69, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b01011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1005,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 69, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b01101000; cin = 1'b1; // Expected: {'sum': 209, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b01101000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1006,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 209, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b10000110; cin = 1'b1; // Expected: {'sum': 67, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b10000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1007,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 67, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b00101111; cin = 1'b0; // Expected: {'sum': 212, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b00101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1008,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 212, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110101; b = 8'b10000010; cin = 1'b1; // Expected: {'sum': 56, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110101; b = 8'b10000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1009,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 56, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b01110000; cin = 1'b0; // Expected: {'sum': 237, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b01110000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1010,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 237, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b10110010; cin = 1'b1; // Expected: {'sum': 187, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b10110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1011,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 187, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b11000101; cin = 1'b1; // Expected: {'sum': 250, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b11000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1012,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 250, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100110; b = 8'b10011110; cin = 1'b1; // Expected: {'sum': 133, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100110; b = 8'b10011110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1013,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 133, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b11110000; cin = 1'b1; // Expected: {'sum': 208, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b11110000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1014,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 208, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b00000100; cin = 1'b1; // Expected: {'sum': 136, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b00000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1015,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 136, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b00011111; cin = 1'b0; // Expected: {'sum': 32, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b00011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1016,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 32, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b11110100; cin = 1'b1; // Expected: {'sum': 140, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b11110100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1017,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 140, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001101; b = 8'b11010010; cin = 1'b0; // Expected: {'sum': 223, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001101; b = 8'b11010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1018,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 223, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b10000100; cin = 1'b1; // Expected: {'sum': 120, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b10000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1019,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 120, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b11101001; cin = 1'b1; // Expected: {'sum': 128, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b11101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1020,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 128, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101011; b = 8'b10010100; cin = 1'b1; // Expected: {'sum': 192, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101011; b = 8'b10010100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1021,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 192, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b00000100; cin = 1'b0; // Expected: {'sum': 164, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b00000100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1022,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 164, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b00001110; cin = 1'b1; // Expected: {'sum': 108, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b00001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1023,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 108, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000000; b = 8'b11001001; cin = 1'b0; // Expected: {'sum': 73, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000000; b = 8'b11001001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1024,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 73, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b01100101; cin = 1'b0; // Expected: {'sum': 97, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b01100101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1025,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 97, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b01010100; cin = 1'b0; // Expected: {'sum': 152, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b01010100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1026,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 152, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b10011110; cin = 1'b0; // Expected: {'sum': 238, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b10011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1027,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 238, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011101; b = 8'b01001000; cin = 1'b1; // Expected: {'sum': 38, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011101; b = 8'b01001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1028,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 38, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b10000010; cin = 1'b1; // Expected: {'sum': 12, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b10000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1029,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110000; b = 8'b10001100; cin = 1'b1; // Expected: {'sum': 253, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110000; b = 8'b10001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1030,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 253, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011010; b = 8'b01101010; cin = 1'b1; // Expected: {'sum': 197, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011010; b = 8'b01101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1031,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 197, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b11000010; cin = 1'b0; // Expected: {'sum': 59, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b11000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1032,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 59, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b11001000; cin = 1'b1; // Expected: {'sum': 231, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b11001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1033,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 231, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b01100100; cin = 1'b0; // Expected: {'sum': 224, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b01100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1034,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 224, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011010; b = 8'b00110010; cin = 1'b1; // Expected: {'sum': 13, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011010; b = 8'b00110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1035,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 13, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b00111010; cin = 1'b0; // Expected: {'sum': 60, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b00111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1036,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 60, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b01000100; cin = 1'b0; // Expected: {'sum': 52, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b01000100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1037,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 52, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b00001001; cin = 1'b1; // Expected: {'sum': 131, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b00001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1038,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 131, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b01111001; cin = 1'b1; // Expected: {'sum': 208, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b01111001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1039,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 208, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011000; b = 8'b10100100; cin = 1'b0; // Expected: {'sum': 252, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011000; b = 8'b10100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1040,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 252, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010110; b = 8'b01110111; cin = 1'b1; // Expected: {'sum': 78, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010110; b = 8'b01110111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1041,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 78, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110011; b = 8'b10001000; cin = 1'b0; // Expected: {'sum': 59, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110011; b = 8'b10001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1042,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 59, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b10011001; cin = 1'b0; // Expected: {'sum': 57, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b10011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1043,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 57, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111101; b = 8'b00001110; cin = 1'b0; // Expected: {'sum': 11, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111101; b = 8'b00001110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1044,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 11, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001100; b = 8'b00100100; cin = 1'b0; // Expected: {'sum': 176, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001100; b = 8'b00100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1045,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 176, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001100; b = 8'b00000011; cin = 1'b0; // Expected: {'sum': 143, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001100; b = 8'b00000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1046,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 143, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b01000000; cin = 1'b1; // Expected: {'sum': 242, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b01000000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1047,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 242, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b10000011; cin = 1'b1; // Expected: {'sum': 200, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b10000011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1048,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 200, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b00100100; cin = 1'b0; // Expected: {'sum': 151, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b00100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1049,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 151, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001110; b = 8'b10110100; cin = 1'b1; // Expected: {'sum': 3, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001110; b = 8'b10110100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1050,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001001; b = 8'b10011011; cin = 1'b0; // Expected: {'sum': 100, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001001; b = 8'b10011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1051,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 100, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000001; b = 8'b01001110; cin = 1'b1; // Expected: {'sum': 16, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000001; b = 8'b01001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1052,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 16, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001100; b = 8'b00010010; cin = 1'b1; // Expected: {'sum': 159, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001100; b = 8'b00010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1053,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 159, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000110; b = 8'b10010011; cin = 1'b1; // Expected: {'sum': 90, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000110; b = 8'b10010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1054,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 90, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b01010000; cin = 1'b1; // Expected: {'sum': 152, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b01010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1055,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 152, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100011; b = 8'b01011010; cin = 1'b1; // Expected: {'sum': 62, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100011; b = 8'b01011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1056,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 62, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110010; b = 8'b01010101; cin = 1'b1; // Expected: {'sum': 200, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110010; b = 8'b01010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1057,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 200, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b01111010; cin = 1'b1; // Expected: {'sum': 216, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b01111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1058,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 216, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b10111111; cin = 1'b1; // Expected: {'sum': 42, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b10111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1059,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 42, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b00001111; cin = 1'b1; // Expected: {'sum': 224, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b00001111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1060,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 224, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000000; b = 8'b01001011; cin = 1'b0; // Expected: {'sum': 203, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000000; b = 8'b01001011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1061,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 203, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b00110001; cin = 1'b0; // Expected: {'sum': 210, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b00110001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1062,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 210, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001001; b = 8'b00110101; cin = 1'b0; // Expected: {'sum': 126, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001001; b = 8'b00110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1063,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 126, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111011; b = 8'b10111001; cin = 1'b0; // Expected: {'sum': 244, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111011; b = 8'b10111001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1064,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 244, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001110; b = 8'b11110010; cin = 1'b0; // Expected: {'sum': 0, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001110; b = 8'b11110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1065,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100111; b = 8'b01011001; cin = 1'b0; // Expected: {'sum': 0, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100111; b = 8'b01011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1066,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b01001101; cin = 1'b0; // Expected: {'sum': 101, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b01001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1067,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 101, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b01000011; cin = 1'b1; // Expected: {'sum': 183, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b01000011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1068,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 183, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b11011111; cin = 1'b1; // Expected: {'sum': 213, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b11011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1069,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 213, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011001; b = 8'b00000110; cin = 1'b0; // Expected: {'sum': 31, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011001; b = 8'b00000110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1070,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 31, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b10001000; cin = 1'b0; // Expected: {'sum': 103, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b10001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1071,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 103, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010100; b = 8'b10111111; cin = 1'b1; // Expected: {'sum': 20, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010100; b = 8'b10111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1072,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 20, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b01010110; cin = 1'b1; // Expected: {'sum': 237, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b01010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1073,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 237, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101111; b = 8'b11001000; cin = 1'b0; // Expected: {'sum': 247, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101111; b = 8'b11001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1074,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 247, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b11001101; cin = 1'b0; // Expected: {'sum': 35, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b11001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1075,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 35, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111000; b = 8'b10010101; cin = 1'b1; // Expected: {'sum': 206, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111000; b = 8'b10010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1076,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 206, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011000; b = 8'b10110111; cin = 1'b0; // Expected: {'sum': 15, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011000; b = 8'b10110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1077,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b00000000; cin = 1'b1; // Expected: {'sum': 109, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b00000000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1078,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 109, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011001; b = 8'b00010000; cin = 1'b1; // Expected: {'sum': 170, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011001; b = 8'b00010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1079,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 170, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b01110101; cin = 1'b0; // Expected: {'sum': 49, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b01110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1080,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 49, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b00011000; cin = 1'b0; // Expected: {'sum': 253, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b00011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1081,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 253, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b00001111; cin = 1'b1; // Expected: {'sum': 153, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b00001111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1082,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 153, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110001; b = 8'b01101101; cin = 1'b1; // Expected: {'sum': 159, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110001; b = 8'b01101101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1083,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 159, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b01100011; cin = 1'b1; // Expected: {'sum': 124, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b01100011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1084,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 124, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b11110111; cin = 1'b0; // Expected: {'sum': 151, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b11110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1085,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 151, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b00011110; cin = 1'b1; // Expected: {'sum': 153, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b00011110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1086,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 153, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b01000111; cin = 1'b1; // Expected: {'sum': 56, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b01000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1087,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 56, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b11011110; cin = 1'b0; // Expected: {'sum': 137, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b11011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1088,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 137, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b01011011; cin = 1'b1; // Expected: {'sum': 46, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b01011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1089,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 46, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b00101100; cin = 1'b1; // Expected: {'sum': 162, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b00101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1090,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 162, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b00010100; cin = 1'b1; // Expected: {'sum': 85, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b00010100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1091,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 85, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b10010001; cin = 1'b0; // Expected: {'sum': 31, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b10010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1092,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 31, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b11010111; cin = 1'b1; // Expected: {'sum': 247, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b11010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1093,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 247, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b11011100; cin = 1'b1; // Expected: {'sum': 89, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b11011100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1094,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 89, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100110; b = 8'b10010101; cin = 1'b1; // Expected: {'sum': 124, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100110; b = 8'b10010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1095,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 124, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000101; b = 8'b10110111; cin = 1'b1; // Expected: {'sum': 125, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000101; b = 8'b10110111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1096,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 125, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011100; b = 8'b01000111; cin = 1'b1; // Expected: {'sum': 36, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011100; b = 8'b01000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1097,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 36, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000011; b = 8'b01001010; cin = 1'b1; // Expected: {'sum': 78, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000011; b = 8'b01001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1098,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 78, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010110; b = 8'b01001000; cin = 1'b0; // Expected: {'sum': 30, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010110; b = 8'b01001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1099,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 30, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b10001110; cin = 1'b0; // Expected: {'sum': 187, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b10001110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1100,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 187, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b11011011; cin = 1'b0; // Expected: {'sum': 143, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b11011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1101,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 143, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001011; b = 8'b00010101; cin = 1'b1; // Expected: {'sum': 97, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001011; b = 8'b00010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1102,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 97, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b01000011; cin = 1'b1; // Expected: {'sum': 177, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b01000011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1103,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 177, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001100; b = 8'b10101101; cin = 1'b0; // Expected: {'sum': 185, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001100; b = 8'b10101101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1104,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 185, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b11100011; cin = 1'b0; // Expected: {'sum': 184, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b11100011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1105,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 184, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b10100101; cin = 1'b0; // Expected: {'sum': 3, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b10100101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1106,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b00001001; cin = 1'b1; // Expected: {'sum': 8, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b00001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1107,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 8, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001100; b = 8'b00011111; cin = 1'b1; // Expected: {'sum': 236, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001100; b = 8'b00011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1108,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 236, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100000; b = 8'b00011011; cin = 1'b1; // Expected: {'sum': 124, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100000; b = 8'b00011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1109,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 124, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b10101110; cin = 1'b1; // Expected: {'sum': 65, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b10101110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1110,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 65, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b00000011; cin = 1'b0; // Expected: {'sum': 186, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b00000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1111,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 186, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100111; b = 8'b11000010; cin = 1'b0; // Expected: {'sum': 41, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100111; b = 8'b11000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1112,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 41, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b01110111; cin = 1'b1; // Expected: {'sum': 13, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b01110111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1113,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 13, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b10100100; cin = 1'b0; // Expected: {'sum': 116, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b10100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1114,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 116, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b01100000; cin = 1'b0; // Expected: {'sum': 203, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b01100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1115,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 203, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b00100001; cin = 1'b0; // Expected: {'sum': 213, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b00100001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1116,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 213, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011110; b = 8'b10000011; cin = 1'b0; // Expected: {'sum': 97, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011110; b = 8'b10000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1117,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 97, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b01110101; cin = 1'b1; // Expected: {'sum': 195, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b01110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1118,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 195, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b01010000; cin = 1'b0; // Expected: {'sum': 53, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b01010000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1119,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 53, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b11101001; cin = 1'b1; // Expected: {'sum': 120, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b11101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1120,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 120, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b11010110; cin = 1'b0; // Expected: {'sum': 12, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b11010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1121,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b01011110; cin = 1'b0; // Expected: {'sum': 95, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b01011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1122,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 95, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b10111000; cin = 1'b0; // Expected: {'sum': 88, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b10111000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1123,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 88, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b10111010; cin = 1'b1; // Expected: {'sum': 2, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b10111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1124,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b01100000; cin = 1'b1; // Expected: {'sum': 197, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b01100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1125,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 197, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b11111010; cin = 1'b0; // Expected: {'sum': 135, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b11111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1126,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 135, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111011; b = 8'b00100000; cin = 1'b0; // Expected: {'sum': 91, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111011; b = 8'b00100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1127,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 91, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b01000110; cin = 1'b0; // Expected: {'sum': 221, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b01000110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1128,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 221, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000110; b = 8'b00111000; cin = 1'b0; // Expected: {'sum': 254, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000110; b = 8'b00111000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1129,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 254, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110100; b = 8'b11000001; cin = 1'b0; // Expected: {'sum': 53, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110100; b = 8'b11000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1130,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 53, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b11001100; cin = 1'b0; // Expected: {'sum': 39, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b11001100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1131,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 39, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101001; b = 8'b10001111; cin = 1'b1; // Expected: {'sum': 121, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101001; b = 8'b10001111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1132,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 121, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001000; b = 8'b00000110; cin = 1'b0; // Expected: {'sum': 206, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001000; b = 8'b00000110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1133,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 206, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011001; b = 8'b10111101; cin = 1'b0; // Expected: {'sum': 22, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011001; b = 8'b10111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1134,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 22, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b01011111; cin = 1'b1; // Expected: {'sum': 203, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b01011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1135,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 203, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b11001110; cin = 1'b1; // Expected: {'sum': 45, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b11001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1136,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 45, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011001; b = 8'b00000111; cin = 1'b1; // Expected: {'sum': 97, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011001; b = 8'b00000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1137,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 97, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011001; b = 8'b00000100; cin = 1'b1; // Expected: {'sum': 94, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011001; b = 8'b00000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1138,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 94, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010001; b = 8'b11110100; cin = 1'b0; // Expected: {'sum': 197, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010001; b = 8'b11110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1139,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 197, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b10000111; cin = 1'b1; // Expected: {'sum': 137, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b10000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1140,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 137, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b00011100; cin = 1'b0; // Expected: {'sum': 132, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b00011100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1141,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 132, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101111; b = 8'b01111100; cin = 1'b1; // Expected: {'sum': 236, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101111; b = 8'b01111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1142,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 236, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b11101110; cin = 1'b1; // Expected: {'sum': 152, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b11101110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1143,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 152, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111010; b = 8'b00110011; cin = 1'b0; // Expected: {'sum': 45, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111010; b = 8'b00110011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1144,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 45, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010101; b = 8'b00001010; cin = 1'b1; // Expected: {'sum': 96, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010101; b = 8'b00001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1145,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 96, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b11000100; cin = 1'b0; // Expected: {'sum': 49, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b11000100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1146,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 49, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b00000011; cin = 1'b0; // Expected: {'sum': 2, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b00000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1147,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011111; b = 8'b11000010; cin = 1'b0; // Expected: {'sum': 33, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011111; b = 8'b11000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1148,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 33, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b11101101; cin = 1'b1; // Expected: {'sum': 239, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b11101101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1149,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 239, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100100; b = 8'b11000100; cin = 1'b1; // Expected: {'sum': 105, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100100; b = 8'b11000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1150,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 105, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b01000010; cin = 1'b0; // Expected: {'sum': 190, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b01000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1151,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 190, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b11001111; cin = 1'b0; // Expected: {'sum': 85, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b11001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1152,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 85, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001110; b = 8'b10100000; cin = 1'b0; // Expected: {'sum': 238, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001110; b = 8'b10100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1153,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 238, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101010; b = 8'b00010010; cin = 1'b1; // Expected: {'sum': 61, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101010; b = 8'b00010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1154,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 61, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b01011110; cin = 1'b1; // Expected: {'sum': 221, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b01011110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1155,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 221, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b00010011; cin = 1'b1; // Expected: {'sum': 149, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b00010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1156,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 149, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b00101110; cin = 1'b1; // Expected: {'sum': 118, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b00101110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1157,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 118, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b11110010; cin = 1'b1; // Expected: {'sum': 21, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b11110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1158,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 21, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b10010111; cin = 1'b0; // Expected: {'sum': 222, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b10010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1159,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 222, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b11100100; cin = 1'b0; // Expected: {'sum': 160, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b11100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1160,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 160, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000011; b = 8'b10010111; cin = 1'b0; // Expected: {'sum': 154, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000011; b = 8'b10010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1161,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 154, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b11000001; cin = 1'b0; // Expected: {'sum': 47, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b11000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1162,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 47, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001111; b = 8'b10011101; cin = 1'b1; // Expected: {'sum': 237, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001111; b = 8'b10011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1163,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 237, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b11110101; cin = 1'b1; // Expected: {'sum': 16, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b11110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1164,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 16, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b10101001; cin = 1'b0; // Expected: {'sum': 174, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b10101001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1165,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 174, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b10011110; cin = 1'b1; // Expected: {'sum': 7, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b10011110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1166,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001011; b = 8'b01101110; cin = 1'b1; // Expected: {'sum': 58, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001011; b = 8'b01101110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1167,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 58, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011011; b = 8'b11100000; cin = 1'b0; // Expected: {'sum': 251, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011011; b = 8'b11100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1168,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 251, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b01010011; cin = 1'b1; // Expected: {'sum': 160, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b01010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1169,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 160, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b00100110; cin = 1'b1; // Expected: {'sum': 103, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b00100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1170,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 103, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111110; b = 8'b10111011; cin = 1'b1; // Expected: {'sum': 250, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111110; b = 8'b10111011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1171,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 250, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b00011010; cin = 1'b0; // Expected: {'sum': 94, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b00011010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1172,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 94, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b00111110; cin = 1'b0; // Expected: {'sum': 189, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b00111110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1173,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 189, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b01011000; cin = 1'b1; // Expected: {'sum': 198, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b01011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1174,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 198, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b10010110; cin = 1'b1; // Expected: {'sum': 75, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b10010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1175,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 75, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b10110110; cin = 1'b1; // Expected: {'sum': 133, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b10110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1176,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 133, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b00101011; cin = 1'b1; // Expected: {'sum': 98, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b00101011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1177,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 98, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000111; b = 8'b11111110; cin = 1'b1; // Expected: {'sum': 134, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000111; b = 8'b11111110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1178,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 134, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b00010100; cin = 1'b1; // Expected: {'sum': 50, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b00010100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1179,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 50, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b10111101; cin = 1'b0; // Expected: {'sum': 48, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b10111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1180,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 48, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b10101001; cin = 1'b1; // Expected: {'sum': 199, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b10101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1181,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 199, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010000; b = 8'b10110001; cin = 1'b0; // Expected: {'sum': 193, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010000; b = 8'b10110001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1182,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 193, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b11010110; cin = 1'b1; // Expected: {'sum': 144, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b11010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1183,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 144, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011101; b = 8'b11010110; cin = 1'b0; // Expected: {'sum': 115, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011101; b = 8'b11010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1184,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 115, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b01111111; cin = 1'b0; // Expected: {'sum': 42, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b01111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1185,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 42, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001000; b = 8'b11111010; cin = 1'b1; // Expected: {'sum': 67, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001000; b = 8'b11111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1186,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 67, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100000; b = 8'b11110010; cin = 1'b1; // Expected: {'sum': 19, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100000; b = 8'b11110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1187,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 19, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b00011101; cin = 1'b1; // Expected: {'sum': 130, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b00011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1188,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 130, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110000; b = 8'b00000000; cin = 1'b1; // Expected: {'sum': 49, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110000; b = 8'b00000000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1189,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 49, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010101; b = 8'b00000010; cin = 1'b0; // Expected: {'sum': 23, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010101; b = 8'b00000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1190,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 23, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010011; b = 8'b01000000; cin = 1'b1; // Expected: {'sum': 148, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010011; b = 8'b01000000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1191,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 148, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b10110111; cin = 1'b0; // Expected: {'sum': 104, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b10110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1192,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 104, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b11011100; cin = 1'b0; // Expected: {'sum': 68, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b11011100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1193,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 68, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b11011110; cin = 1'b1; // Expected: {'sum': 108, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b11011110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1194,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 108, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b00010001; cin = 1'b1; // Expected: {'sum': 140, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b00010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1195,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 140, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b01010000; cin = 1'b0; // Expected: {'sum': 255, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b01010000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1196,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 255, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b00011100; cin = 1'b1; // Expected: {'sum': 105, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b00011100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1197,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 105, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101110; b = 8'b01011010; cin = 1'b1; // Expected: {'sum': 137, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101110; b = 8'b01011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1198,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 137, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011001; b = 8'b11101000; cin = 1'b0; // Expected: {'sum': 65, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011001; b = 8'b11101000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1199,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 65, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b10000010; cin = 1'b0; // Expected: {'sum': 138, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b10000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1200,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 138, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b10001000; cin = 1'b1; // Expected: {'sum': 252, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b10001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1201,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 252, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001001; b = 8'b10111000; cin = 1'b1; // Expected: {'sum': 2, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001001; b = 8'b10111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1202,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b01000001; cin = 1'b1; // Expected: {'sum': 83, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b01000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1203,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 83, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b10000000; cin = 1'b1; // Expected: {'sum': 122, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b10000000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1204,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 122, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b01010011; cin = 1'b0; // Expected: {'sum': 227, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b01010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1205,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 227, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b00010001; cin = 1'b1; // Expected: {'sum': 208, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b00010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1206,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 208, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b00010100; cin = 1'b0; // Expected: {'sum': 94, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b00010100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1207,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 94, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b11101111; cin = 1'b0; // Expected: {'sum': 41, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b11101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1208,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 41, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011010; b = 8'b10100110; cin = 1'b1; // Expected: {'sum': 129, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011010; b = 8'b10100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1209,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 129, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000000; b = 8'b00001100; cin = 1'b0; // Expected: {'sum': 140, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000000; b = 8'b00001100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1210,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 140, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b11000011; cin = 1'b0; // Expected: {'sum': 13, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b11000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1211,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 13, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b11010010; cin = 1'b1; // Expected: {'sum': 132, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b11010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1212,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 132, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b10111000; cin = 1'b1; // Expected: {'sum': 90, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b10111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1213,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 90, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b11010010; cin = 1'b1; // Expected: {'sum': 75, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b11010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1214,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 75, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b01110111; cin = 1'b0; // Expected: {'sum': 34, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b01110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1215,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 34, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b00111011; cin = 1'b0; // Expected: {'sum': 22, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b00111011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1216,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 22, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b01000001; cin = 1'b0; // Expected: {'sum': 220, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b01000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1217,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 220, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b00010011; cin = 1'b0; // Expected: {'sum': 0, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b00010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1218,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b00100111; cin = 1'b0; // Expected: {'sum': 158, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b00100111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1219,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 158, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b01011111; cin = 1'b1; // Expected: {'sum': 247, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b01011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1220,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 247, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111110; b = 8'b00011010; cin = 1'b1; // Expected: {'sum': 89, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111110; b = 8'b00011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1221,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 89, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b11010011; cin = 1'b0; // Expected: {'sum': 64, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b11010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1222,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 64, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b00111011; cin = 1'b1; // Expected: {'sum': 235, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b00111011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1223,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 235, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110101; b = 8'b00101010; cin = 1'b0; // Expected: {'sum': 95, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110101; b = 8'b00101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1224,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 95, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b10001001; cin = 1'b1; // Expected: {'sum': 98, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b10001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1225,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 98, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b00100100; cin = 1'b1; // Expected: {'sum': 167, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b00100100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1226,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 167, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b10100001; cin = 1'b0; // Expected: {'sum': 146, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b10100001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1227,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 146, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b00010101; cin = 1'b1; // Expected: {'sum': 132, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b00010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1228,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 132, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b01111001; cin = 1'b1; // Expected: {'sum': 156, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b01111001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1229,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 156, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100111; b = 8'b00000000; cin = 1'b0; // Expected: {'sum': 231, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100111; b = 8'b00000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1230,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 231, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000110; b = 8'b00011110; cin = 1'b0; // Expected: {'sum': 228, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000110; b = 8'b00011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1231,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 228, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b10100110; cin = 1'b1; // Expected: {'sum': 19, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b10100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1232,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 19, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b01110011; cin = 1'b1; // Expected: {'sum': 248, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b01110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1233,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 248, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b10100101; cin = 1'b1; // Expected: {'sum': 56, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b10100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1234,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 56, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001111; b = 8'b11100000; cin = 1'b1; // Expected: {'sum': 48, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001111; b = 8'b11100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1235,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 48, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b01011111; cin = 1'b1; // Expected: {'sum': 75, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b01011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1236,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 75, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100111; b = 8'b10110000; cin = 1'b1; // Expected: {'sum': 88, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100111; b = 8'b10110000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1237,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 88, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101101; b = 8'b01101001; cin = 1'b1; // Expected: {'sum': 23, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101101; b = 8'b01101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1238,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 23, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b01000111; cin = 1'b1; // Expected: {'sum': 73, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b01000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1239,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 73, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100000; b = 8'b10100111; cin = 1'b0; // Expected: {'sum': 7, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100000; b = 8'b10100111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1240,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b11110001; cin = 1'b0; // Expected: {'sum': 86, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b11110001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1241,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 86, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011101; b = 8'b10100000; cin = 1'b0; // Expected: {'sum': 125, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011101; b = 8'b10100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1242,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 125, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010101; b = 8'b01111111; cin = 1'b1; // Expected: {'sum': 149, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010101; b = 8'b01111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1243,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 149, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b00001111; cin = 1'b0; // Expected: {'sum': 116, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b00001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1244,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 116, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b11000111; cin = 1'b1; // Expected: {'sum': 169, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b11000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1245,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 169, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b01010111; cin = 1'b0; // Expected: {'sum': 47, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b01010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1246,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 47, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b11010101; cin = 1'b0; // Expected: {'sum': 94, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b11010101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1247,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 94, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110001; b = 8'b01001110; cin = 1'b0; // Expected: {'sum': 191, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110001; b = 8'b01001110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1248,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 191, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b01010001; cin = 1'b1; // Expected: {'sum': 188, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b01010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1249,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 188, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100000; b = 8'b10001100; cin = 1'b1; // Expected: {'sum': 173, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100000; b = 8'b10001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1250,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 173, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b00010111; cin = 1'b0; // Expected: {'sum': 89, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b00010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1251,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 89, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100011; b = 8'b00110001; cin = 1'b1; // Expected: {'sum': 21, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100011; b = 8'b00110001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1252,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 21, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b00011000; cin = 1'b0; // Expected: {'sum': 60, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b00011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1253,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 60, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b10011101; cin = 1'b0; // Expected: {'sum': 42, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b10011101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1254,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 42, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b10110010; cin = 1'b1; // Expected: {'sum': 92, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b10110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1255,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 92, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110010; b = 8'b11010111; cin = 1'b0; // Expected: {'sum': 73, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110010; b = 8'b11010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1256,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 73, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b10101011; cin = 1'b1; // Expected: {'sum': 198, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b10101011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1257,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 198, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b11010110; cin = 1'b1; // Expected: {'sum': 103, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b11010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1258,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 103, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b11011100; cin = 1'b1; // Expected: {'sum': 59, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b11011100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1259,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 59, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011010; b = 8'b10001010; cin = 1'b1; // Expected: {'sum': 101, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011010; b = 8'b10001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1260,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 101, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b01011011; cin = 1'b1; // Expected: {'sum': 68, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b01011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1261,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 68, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b00001000; cin = 1'b1; // Expected: {'sum': 155, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b00001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1262,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 155, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b00000110; cin = 1'b1; // Expected: {'sum': 199, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b00000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1263,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 199, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b01100010; cin = 1'b0; // Expected: {'sum': 152, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b01100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1264,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 152, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010001; b = 8'b01010110; cin = 1'b1; // Expected: {'sum': 40, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010001; b = 8'b01010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1265,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 40, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b10001111; cin = 1'b1; // Expected: {'sum': 131, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b10001111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1266,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 131, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b11101111; cin = 1'b1; // Expected: {'sum': 60, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b11101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1267,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 60, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010100; b = 8'b01010010; cin = 1'b0; // Expected: {'sum': 102, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010100; b = 8'b01010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1268,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 102, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b01111101; cin = 1'b0; // Expected: {'sum': 15, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b01111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1269,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101100; b = 8'b00100110; cin = 1'b1; // Expected: {'sum': 19, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101100; b = 8'b00100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1270,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 19, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b11011001; cin = 1'b1; // Expected: {'sum': 206, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b11011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1271,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 206, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b00101010; cin = 1'b0; // Expected: {'sum': 134, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b00101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1272,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 134, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100000; b = 8'b10010010; cin = 1'b0; // Expected: {'sum': 178, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100000; b = 8'b10010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1273,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 178, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b11111011; cin = 1'b0; // Expected: {'sum': 137, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b11111011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1274,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 137, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b00001100; cin = 1'b1; // Expected: {'sum': 117, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b00001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1275,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 117, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000011; b = 8'b00111110; cin = 1'b1; // Expected: {'sum': 2, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000011; b = 8'b00111110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1276,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001000; b = 8'b10010001; cin = 1'b1; // Expected: {'sum': 90, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001000; b = 8'b10010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1277,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 90, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b01000101; cin = 1'b1; // Expected: {'sum': 60, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b01000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1278,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 60, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b11101100; cin = 1'b1; // Expected: {'sum': 187, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b11101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1279,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 187, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111001; b = 8'b10100000; cin = 1'b1; // Expected: {'sum': 218, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111001; b = 8'b10100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1280,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 218, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b10001101; cin = 1'b1; // Expected: {'sum': 161, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b10001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1281,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 161, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101101; b = 8'b11011001; cin = 1'b0; // Expected: {'sum': 134, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101101; b = 8'b11011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1282,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 134, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b11100100; cin = 1'b1; // Expected: {'sum': 139, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b11100100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1283,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 139, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010011; b = 8'b00111111; cin = 1'b1; // Expected: {'sum': 19, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010011; b = 8'b00111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1284,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 19, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111011; b = 8'b10100000; cin = 1'b1; // Expected: {'sum': 28, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111011; b = 8'b10100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1285,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 28, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111011; b = 8'b10010011; cin = 1'b0; // Expected: {'sum': 206, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111011; b = 8'b10010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1286,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 206, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100000; b = 8'b01101101; cin = 1'b0; // Expected: {'sum': 77, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100000; b = 8'b01101101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1287,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 77, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b10010101; cin = 1'b1; // Expected: {'sum': 179, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b10010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1288,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 179, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011111; b = 8'b11011011; cin = 1'b0; // Expected: {'sum': 122, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011111; b = 8'b11011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1289,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 122, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000110; b = 8'b00001110; cin = 1'b1; // Expected: {'sum': 85, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000110; b = 8'b00001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1290,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 85, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b11011111; cin = 1'b1; // Expected: {'sum': 9, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b11011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1291,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 9, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b01111010; cin = 1'b0; // Expected: {'sum': 5, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b01111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1292,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 5, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b11100110; cin = 1'b1; // Expected: {'sum': 161, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b11100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1293,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 161, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110010; b = 8'b00010100; cin = 1'b0; // Expected: {'sum': 134, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110010; b = 8'b00010100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1294,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 134, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b11110101; cin = 1'b0; // Expected: {'sum': 250, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b11110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1295,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 250, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b00101001; cin = 1'b1; // Expected: {'sum': 171, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b00101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1296,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 171, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000101; b = 8'b00011001; cin = 1'b0; // Expected: {'sum': 158, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000101; b = 8'b00011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1297,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 158, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001010; b = 8'b00110100; cin = 1'b0; // Expected: {'sum': 190, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001010; b = 8'b00110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1298,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 190, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000011; b = 8'b00111010; cin = 1'b0; // Expected: {'sum': 61, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000011; b = 8'b00111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1299,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 61, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101001; b = 8'b00010111; cin = 1'b1; // Expected: {'sum': 1, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101001; b = 8'b00010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1300,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b11001111; cin = 1'b1; // Expected: {'sum': 239, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b11001111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1301,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 239, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100000; b = 8'b11010011; cin = 1'b1; // Expected: {'sum': 52, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100000; b = 8'b11010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1302,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 52, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100000; b = 8'b10110010; cin = 1'b1; // Expected: {'sum': 147, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100000; b = 8'b10110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1303,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 147, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011110; b = 8'b00101101; cin = 1'b1; // Expected: {'sum': 12, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011110; b = 8'b00101101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1304,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b00011100; cin = 1'b0; // Expected: {'sum': 179, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b00011100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1305,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 179, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b10011000; cin = 1'b1; // Expected: {'sum': 221, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b10011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1306,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 221, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b11101111; cin = 1'b0; // Expected: {'sum': 220, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b11101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1307,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 220, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b11111101; cin = 1'b0; // Expected: {'sum': 95, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b11111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1308,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 95, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000111; b = 8'b01111110; cin = 1'b1; // Expected: {'sum': 70, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000111; b = 8'b01111110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1309,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 70, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111000; b = 8'b01010011; cin = 1'b0; // Expected: {'sum': 75, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111000; b = 8'b01010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1310,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 75, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010011; b = 8'b00100110; cin = 1'b0; // Expected: {'sum': 185, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010011; b = 8'b00100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1311,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 185, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b11001010; cin = 1'b1; // Expected: {'sum': 5, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b11001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1312,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 5, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000001; b = 8'b10010110; cin = 1'b1; // Expected: {'sum': 88, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000001; b = 8'b10010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1313,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 88, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000011; b = 8'b11011110; cin = 1'b0; // Expected: {'sum': 225, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000011; b = 8'b11011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1314,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 225, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b11110010; cin = 1'b1; // Expected: {'sum': 94, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b11110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1315,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 94, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001011; b = 8'b00011010; cin = 1'b0; // Expected: {'sum': 37, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001011; b = 8'b00011010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1316,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 37, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b11010010; cin = 1'b1; // Expected: {'sum': 149, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b11010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1317,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 149, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b01000001; cin = 1'b0; // Expected: {'sum': 22, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b01000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1318,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 22, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110001; b = 8'b10110101; cin = 1'b1; // Expected: {'sum': 39, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110001; b = 8'b10110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1319,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 39, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b01110011; cin = 1'b1; // Expected: {'sum': 118, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b01110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1320,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 118, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b01101010; cin = 1'b0; // Expected: {'sum': 147, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b01101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1321,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 147, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b01000111; cin = 1'b0; // Expected: {'sum': 59, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b01000111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1322,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 59, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000111; b = 8'b01001111; cin = 1'b0; // Expected: {'sum': 22, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000111; b = 8'b01001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1323,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 22, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b01011000; cin = 1'b1; // Expected: {'sum': 169, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b01011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1324,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 169, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111101; b = 8'b10101001; cin = 1'b0; // Expected: {'sum': 166, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111101; b = 8'b10101001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1325,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 166, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b11110010; cin = 1'b0; // Expected: {'sum': 252, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b11110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1326,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 252, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b10011011; cin = 1'b1; // Expected: {'sum': 117, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b10011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1327,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 117, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b00001111; cin = 1'b0; // Expected: {'sum': 192, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b00001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1328,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 192, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b10101101; cin = 1'b0; // Expected: {'sum': 53, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b10101101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1329,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 53, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100111; b = 8'b10110101; cin = 1'b1; // Expected: {'sum': 157, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100111; b = 8'b10110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1330,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 157, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b01101000; cin = 1'b1; // Expected: {'sum': 244, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b01101000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1331,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 244, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010101; b = 8'b00010100; cin = 1'b0; // Expected: {'sum': 105, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010101; b = 8'b00010100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1332,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 105, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100111; b = 8'b10001111; cin = 1'b0; // Expected: {'sum': 182, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100111; b = 8'b10001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1333,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 182, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b10001111; cin = 1'b0; // Expected: {'sum': 4, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b10001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1334,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000110; b = 8'b01011110; cin = 1'b1; // Expected: {'sum': 165, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000110; b = 8'b01011110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1335,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 165, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b11100001; cin = 1'b1; // Expected: {'sum': 0, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b11100001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1336,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b00110101; cin = 1'b1; // Expected: {'sum': 217, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b00110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1337,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 217, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b01100000; cin = 1'b0; // Expected: {'sum': 80, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b01100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1338,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 80, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b10100010; cin = 1'b1; // Expected: {'sum': 163, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b10100010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1339,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 163, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b01011001; cin = 1'b1; // Expected: {'sum': 190, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b01011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1340,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 190, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110101; b = 8'b11111111; cin = 1'b1; // Expected: {'sum': 53, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110101; b = 8'b11111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1341,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 53, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b11000001; cin = 1'b1; // Expected: {'sum': 144, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b11000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1342,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 144, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b01011111; cin = 1'b0; // Expected: {'sum': 24, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b01011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1343,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 24, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011010; b = 8'b10010011; cin = 1'b1; // Expected: {'sum': 110, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011010; b = 8'b10010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1344,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 110, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b10010111; cin = 1'b0; // Expected: {'sum': 64, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b10010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1345,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 64, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110111; b = 8'b10101100; cin = 1'b0; // Expected: {'sum': 227, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110111; b = 8'b10101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1346,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 227, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b11001010; cin = 1'b1; // Expected: {'sum': 238, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b11001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1347,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 238, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101100; b = 8'b10101000; cin = 1'b1; // Expected: {'sum': 85, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101100; b = 8'b10101000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1348,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 85, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b01011110; cin = 1'b1; // Expected: {'sum': 35, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b01011110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1349,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 35, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011011; b = 8'b01010101; cin = 1'b0; // Expected: {'sum': 112, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011011; b = 8'b01010101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1350,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 112, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b00001001; cin = 1'b0; // Expected: {'sum': 83, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b00001001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1351,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 83, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b10111101; cin = 1'b0; // Expected: {'sum': 121, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b10111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1352,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 121, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b01111110; cin = 1'b1; // Expected: {'sum': 213, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b01111110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1353,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 213, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b00001101; cin = 1'b0; // Expected: {'sum': 199, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b00001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1354,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 199, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b10101001; cin = 1'b1; // Expected: {'sum': 157, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b10101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1355,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 157, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011110; b = 8'b01010010; cin = 1'b1; // Expected: {'sum': 49, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011110; b = 8'b01010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1356,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 49, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000110; b = 8'b11101101; cin = 1'b0; // Expected: {'sum': 243, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000110; b = 8'b11101101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1357,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 243, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b00101101; cin = 1'b0; // Expected: {'sum': 247, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b00101101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1358,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 247, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000001; b = 8'b00011010; cin = 1'b1; // Expected: {'sum': 220, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000001; b = 8'b00011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1359,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 220, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b00101110; cin = 1'b0; // Expected: {'sum': 155, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b00101110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1360,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 155, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011111; b = 8'b10111111; cin = 1'b0; // Expected: {'sum': 94, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011111; b = 8'b10111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1361,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 94, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b11110111; cin = 1'b1; // Expected: {'sum': 188, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b11110111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1362,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 188, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110110; b = 8'b11100001; cin = 1'b1; // Expected: {'sum': 88, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110110; b = 8'b11100001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1363,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 88, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b11001010; cin = 1'b1; // Expected: {'sum': 182, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b11001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1364,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 182, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101010; b = 8'b11000110; cin = 1'b1; // Expected: {'sum': 241, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101010; b = 8'b11000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1365,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 241, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000111; b = 8'b11110011; cin = 1'b1; // Expected: {'sum': 123, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000111; b = 8'b11110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1366,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 123, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b11011011; cin = 1'b1; // Expected: {'sum': 132, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b11011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1367,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 132, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100110; b = 8'b00001010; cin = 1'b0; // Expected: {'sum': 48, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100110; b = 8'b00001010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1368,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 48, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b10010101; cin = 1'b0; // Expected: {'sum': 15, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b10010101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1369,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b10011011; cin = 1'b1; // Expected: {'sum': 224, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b10011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1370,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 224, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010101; b = 8'b10000100; cin = 1'b1; // Expected: {'sum': 154, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010101; b = 8'b10000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1371,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 154, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001100; b = 8'b00111010; cin = 1'b1; // Expected: {'sum': 7, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001100; b = 8'b00111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1372,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111101; b = 8'b01101110; cin = 1'b1; // Expected: {'sum': 108, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111101; b = 8'b01101110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1373,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 108, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b10111010; cin = 1'b0; // Expected: {'sum': 149, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b10111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1374,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 149, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b11110001; cin = 1'b0; // Expected: {'sum': 202, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b11110001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1375,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 202, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b00010001; cin = 1'b0; // Expected: {'sum': 211, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b00010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1376,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 211, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110111; b = 8'b11110000; cin = 1'b0; // Expected: {'sum': 39, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110111; b = 8'b11110000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1377,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 39, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b11011000; cin = 1'b0; // Expected: {'sum': 140, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b11011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1378,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 140, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b00110101; cin = 1'b1; // Expected: {'sum': 145, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b00110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1379,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 145, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110001; b = 8'b11011111; cin = 1'b1; // Expected: {'sum': 17, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110001; b = 8'b11011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1380,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 17, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b11011110; cin = 1'b0; // Expected: {'sum': 213, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b11011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1381,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 213, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b11001010; cin = 1'b1; // Expected: {'sum': 162, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b11001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1382,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 162, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b10011100; cin = 1'b1; // Expected: {'sum': 118, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b10011100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1383,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 118, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b01100111; cin = 1'b1; // Expected: {'sum': 230, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b01100111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1384,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 230, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b01100100; cin = 1'b1; // Expected: {'sum': 1, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b01100100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1385,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b11001100; cin = 1'b1; // Expected: {'sum': 9, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b11001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1386,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 9, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b11111101; cin = 1'b0; // Expected: {'sum': 119, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b11111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1387,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 119, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111011; b = 8'b01010111; cin = 1'b1; // Expected: {'sum': 211, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111011; b = 8'b01010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1388,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 211, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b11111000; cin = 1'b1; // Expected: {'sum': 218, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b11111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1389,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 218, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b01010001; cin = 1'b0; // Expected: {'sum': 131, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b01010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1390,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 131, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101010; b = 8'b01110010; cin = 1'b0; // Expected: {'sum': 28, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101010; b = 8'b01110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1391,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 28, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b01011001; cin = 1'b1; // Expected: {'sum': 131, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b01011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1392,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 131, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b01000000; cin = 1'b0; // Expected: {'sum': 150, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b01000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1393,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 150, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b11111000; cin = 1'b0; // Expected: {'sum': 90, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b11111000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1394,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 90, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001110; b = 8'b01110110; cin = 1'b1; // Expected: {'sum': 133, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001110; b = 8'b01110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1395,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 133, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b10001010; cin = 1'b0; // Expected: {'sum': 190, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b10001010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1396,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 190, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010011; b = 8'b01110101; cin = 1'b1; // Expected: {'sum': 9, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010011; b = 8'b01110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1397,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 9, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b10000110; cin = 1'b0; // Expected: {'sum': 8, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b10000110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1398,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 8, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b01100001; cin = 1'b0; // Expected: {'sum': 17, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b01100001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1399,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 17, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010010; b = 8'b10111111; cin = 1'b1; // Expected: {'sum': 210, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010010; b = 8'b10111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1400,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 210, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101111; b = 8'b00101110; cin = 1'b0; // Expected: {'sum': 157, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101111; b = 8'b00101110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1401,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 157, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b01110100; cin = 1'b1; // Expected: {'sum': 171, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b01110100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1402,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 171, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100000; b = 8'b01000110; cin = 1'b1; // Expected: {'sum': 39, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100000; b = 8'b01000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1403,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 39, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b01000110; cin = 1'b1; // Expected: {'sum': 227, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b01000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1404,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 227, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b00010001; cin = 1'b1; // Expected: {'sum': 117, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b00010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1405,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 117, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b10101001; cin = 1'b1; // Expected: {'sum': 146, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b10101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1406,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 146, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b00011110; cin = 1'b0; // Expected: {'sum': 172, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b00011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1407,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 172, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b01101100; cin = 1'b1; // Expected: {'sum': 29, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b01101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1408,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 29, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b00101011; cin = 1'b1; // Expected: {'sum': 240, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b00101011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1409,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 240, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100111; b = 8'b01111100; cin = 1'b1; // Expected: {'sum': 164, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100111; b = 8'b01111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1410,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 164, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b10000000; cin = 1'b0; // Expected: {'sum': 66, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b10000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1411,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 66, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b10011010; cin = 1'b1; // Expected: {'sum': 0, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b10011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1412,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b10110001; cin = 1'b0; // Expected: {'sum': 196, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b10110001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1413,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 196, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101001; b = 8'b10000100; cin = 1'b1; // Expected: {'sum': 110, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101001; b = 8'b10000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1414,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 110, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b01010111; cin = 1'b0; // Expected: {'sum': 95, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b01010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1415,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 95, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101111; b = 8'b00110011; cin = 1'b0; // Expected: {'sum': 34, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101111; b = 8'b00110011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1416,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 34, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010001; b = 8'b01110010; cin = 1'b1; // Expected: {'sum': 68, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010001; b = 8'b01110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1417,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 68, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011010; b = 8'b01101000; cin = 1'b0; // Expected: {'sum': 66, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011010; b = 8'b01101000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1418,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 66, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b10101001; cin = 1'b1; // Expected: {'sum': 130, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b10101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1419,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 130, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111000; b = 8'b01001111; cin = 1'b0; // Expected: {'sum': 71, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111000; b = 8'b01001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1420,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 71, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b01110111; cin = 1'b1; // Expected: {'sum': 40, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b01110111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1421,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 40, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010011; b = 8'b11010001; cin = 1'b0; // Expected: {'sum': 36, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010011; b = 8'b11010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1422,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 36, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010100; b = 8'b11011011; cin = 1'b0; // Expected: {'sum': 47, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010100; b = 8'b11011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1423,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 47, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b10111100; cin = 1'b0; // Expected: {'sum': 124, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b10111100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1424,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 124, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b01011000; cin = 1'b1; // Expected: {'sum': 113, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b01011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1425,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 113, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b11100110; cin = 1'b1; // Expected: {'sum': 250, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b11100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1426,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 250, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b01101010; cin = 1'b0; // Expected: {'sum': 252, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b01101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1427,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 252, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b00100101; cin = 1'b1; // Expected: {'sum': 193, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b00100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1428,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 193, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b00100110; cin = 1'b0; // Expected: {'sum': 129, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b00100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1429,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 129, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100111; b = 8'b00011101; cin = 1'b0; // Expected: {'sum': 196, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100111; b = 8'b00011101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1430,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 196, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000101; b = 8'b10011111; cin = 1'b1; // Expected: {'sum': 101, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000101; b = 8'b10011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1431,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 101, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b01000111; cin = 1'b0; // Expected: {'sum': 52, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b01000111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1432,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 52, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b10100010; cin = 1'b1; // Expected: {'sum': 84, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b10100010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1433,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 84, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b00100000; cin = 1'b0; // Expected: {'sum': 159, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b00100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1434,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 159, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b10100001; cin = 1'b1; // Expected: {'sum': 179, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b10100001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1435,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 179, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110101; b = 8'b11101100; cin = 1'b1; // Expected: {'sum': 34, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110101; b = 8'b11101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1436,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 34, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b10111001; cin = 1'b0; // Expected: {'sum': 230, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b10111001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1437,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 230, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010100; b = 8'b11011111; cin = 1'b0; // Expected: {'sum': 51, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010100; b = 8'b11011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1438,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 51, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b01001001; cin = 1'b1; // Expected: {'sum': 82, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b01001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1439,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 82, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b01011110; cin = 1'b1; // Expected: {'sum': 126, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b01011110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1440,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 126, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b10010001; cin = 1'b1; // Expected: {'sum': 20, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b10010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1441,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 20, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b00100111; cin = 1'b1; // Expected: {'sum': 0, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b00100111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1442,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b10000000; cin = 1'b0; // Expected: {'sum': 208, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b10000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1443,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 208, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b10110110; cin = 1'b1; // Expected: {'sum': 233, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b10110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1444,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 233, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b00000011; cin = 1'b0; // Expected: {'sum': 191, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b00000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1445,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 191, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b00011011; cin = 1'b1; // Expected: {'sum': 169, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b00011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1446,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 169, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111000; b = 8'b00011011; cin = 1'b1; // Expected: {'sum': 84, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111000; b = 8'b00011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1447,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 84, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b01100011; cin = 1'b0; // Expected: {'sum': 175, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b01100011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1448,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 175, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111110; b = 8'b11011010; cin = 1'b0; // Expected: {'sum': 24, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111110; b = 8'b11011010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1449,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 24, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b10111000; cin = 1'b1; // Expected: {'sum': 121, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b10111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1450,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 121, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b11100100; cin = 1'b0; // Expected: {'sum': 251, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b11100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1451,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 251, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101010; b = 8'b01110000; cin = 1'b1; // Expected: {'sum': 91, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101010; b = 8'b01110000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1452,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 91, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b10110110; cin = 1'b1; // Expected: {'sum': 192, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b10110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1453,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 192, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100111; b = 8'b00010011; cin = 1'b1; // Expected: {'sum': 187, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100111; b = 8'b00010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1454,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 187, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101100; b = 8'b01011110; cin = 1'b0; // Expected: {'sum': 10, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101100; b = 8'b01011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1455,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100110; b = 8'b11001000; cin = 1'b0; // Expected: {'sum': 238, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100110; b = 8'b11001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1456,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 238, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010010; b = 8'b01110101; cin = 1'b1; // Expected: {'sum': 136, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010010; b = 8'b01110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1457,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 136, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b10011010; cin = 1'b1; // Expected: {'sum': 76, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b10011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1458,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 76, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b00011101; cin = 1'b0; // Expected: {'sum': 36, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b00011101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1459,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 36, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b00000101; cin = 1'b1; // Expected: {'sum': 184, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b00000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1460,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 184, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010011; b = 8'b01100111; cin = 1'b0; // Expected: {'sum': 186, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010011; b = 8'b01100111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1461,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 186, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b00110101; cin = 1'b1; // Expected: {'sum': 43, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b00110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1462,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 43, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b11101010; cin = 1'b1; // Expected: {'sum': 45, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b11101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1463,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 45, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b01100010; cin = 1'b1; // Expected: {'sum': 62, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b01100010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1464,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 62, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b10000101; cin = 1'b1; // Expected: {'sum': 226, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b10000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1465,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 226, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100111; b = 8'b11001110; cin = 1'b0; // Expected: {'sum': 181, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100111; b = 8'b11001110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1466,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 181, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b11010110; cin = 1'b0; // Expected: {'sum': 134, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b11010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1467,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 134, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b10110011; cin = 1'b0; // Expected: {'sum': 169, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b10110011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1468,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 169, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001110; b = 8'b11110001; cin = 1'b0; // Expected: {'sum': 255, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001110; b = 8'b11110001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1469,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 255, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011110; b = 8'b00100010; cin = 1'b1; // Expected: {'sum': 1, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011110; b = 8'b00100010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1470,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b10100101; cin = 1'b1; // Expected: {'sum': 194, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b10100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1471,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 194, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100110; b = 8'b10111100; cin = 1'b0; // Expected: {'sum': 226, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100110; b = 8'b10111100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1472,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 226, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b00110001; cin = 1'b1; // Expected: {'sum': 22, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b00110001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1473,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 22, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011010; b = 8'b01110011; cin = 1'b1; // Expected: {'sum': 78, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011010; b = 8'b01110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1474,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 78, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111001; b = 8'b01110111; cin = 1'b0; // Expected: {'sum': 176, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111001; b = 8'b01110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1475,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 176, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b00001001; cin = 1'b1; // Expected: {'sum': 194, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b00001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1476,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 194, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100111; b = 8'b11111110; cin = 1'b0; // Expected: {'sum': 229, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100111; b = 8'b11111110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1477,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 229, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101110; b = 8'b01000001; cin = 1'b1; // Expected: {'sum': 112, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101110; b = 8'b01000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1478,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 112, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b11100000; cin = 1'b0; // Expected: {'sum': 19, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b11100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1479,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 19, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b11000000; cin = 1'b0; // Expected: {'sum': 201, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b11000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1480,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 201, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b10100101; cin = 1'b1; // Expected: {'sum': 246, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b10100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1481,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 246, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b11000010; cin = 1'b0; // Expected: {'sum': 48, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b11000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1482,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 48, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100011; b = 8'b11000101; cin = 1'b1; // Expected: {'sum': 169, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100011; b = 8'b11000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1483,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 169, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b00111101; cin = 1'b0; // Expected: {'sum': 243, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b00111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1484,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 243, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010110; b = 8'b11000000; cin = 1'b0; // Expected: {'sum': 150, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010110; b = 8'b11000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1485,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 150, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b01011100; cin = 1'b1; // Expected: {'sum': 3, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b01011100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1486,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b00010110; cin = 1'b1; // Expected: {'sum': 166, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b00010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1487,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 166, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b00100110; cin = 1'b1; // Expected: {'sum': 138, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b00100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1488,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 138, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110100; b = 8'b10000010; cin = 1'b1; // Expected: {'sum': 247, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110100; b = 8'b10000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1489,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 247, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b00101010; cin = 1'b1; // Expected: {'sum': 36, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b00101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1490,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 36, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b11000101; cin = 1'b1; // Expected: {'sum': 102, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b11000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1491,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 102, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b11011101; cin = 1'b0; // Expected: {'sum': 221, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b11011101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1492,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 221, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b01110001; cin = 1'b1; // Expected: {'sum': 205, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b01110001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1493,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 205, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111111; b = 8'b00110011; cin = 1'b0; // Expected: {'sum': 114, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111111; b = 8'b00110011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1494,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 114, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b01010101; cin = 1'b0; // Expected: {'sum': 245, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b01010101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1495,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 245, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001010; b = 8'b10001101; cin = 1'b1; // Expected: {'sum': 24, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001010; b = 8'b10001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1496,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 24, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b10110101; cin = 1'b1; // Expected: {'sum': 60, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b10110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1497,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 60, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b10010100; cin = 1'b1; // Expected: {'sum': 241, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b10010100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1498,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 241, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000100; b = 8'b11011111; cin = 1'b0; // Expected: {'sum': 227, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000100; b = 8'b11011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1499,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 227, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b11111100; cin = 1'b1; // Expected: {'sum': 112, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b11111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1500,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 112, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b00100110; cin = 1'b0; // Expected: {'sum': 11, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b00100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1501,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 11, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b01100000; cin = 1'b1; // Expected: {'sum': 57, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b01100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1502,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 57, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b11011100; cin = 1'b1; // Expected: {'sum': 136, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b11011100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1503,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 136, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b10101011; cin = 1'b0; // Expected: {'sum': 188, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b10101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1504,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 188, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011111; b = 8'b10110100; cin = 1'b1; // Expected: {'sum': 84, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011111; b = 8'b10110100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1505,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 84, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b01000000; cin = 1'b1; // Expected: {'sum': 25, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b01000000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1506,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 25, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b01111111; cin = 1'b1; // Expected: {'sum': 205, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b01111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1507,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 205, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b01000111; cin = 1'b0; // Expected: {'sum': 205, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b01000111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1508,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 205, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b01111001; cin = 1'b1; // Expected: {'sum': 141, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b01111001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1509,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 141, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b01110000; cin = 1'b0; // Expected: {'sum': 91, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b01110000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1510,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 91, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100110; b = 8'b00001110; cin = 1'b1; // Expected: {'sum': 117, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100110; b = 8'b00001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1511,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 117, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b10011001; cin = 1'b0; // Expected: {'sum': 58, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b10011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1512,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 58, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b01110111; cin = 1'b0; // Expected: {'sum': 47, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b01110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1513,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 47, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b10001111; cin = 1'b1; // Expected: {'sum': 194, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b10001111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1514,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 194, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b01110011; cin = 1'b1; // Expected: {'sum': 123, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b01110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1515,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 123, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b10011100; cin = 1'b0; // Expected: {'sum': 138, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b10011100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1516,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 138, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b10111001; cin = 1'b1; // Expected: {'sum': 168, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b10111001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1517,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 168, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b00010111; cin = 1'b1; // Expected: {'sum': 98, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b00010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1518,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 98, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b11110010; cin = 1'b1; // Expected: {'sum': 123, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b11110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1519,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 123, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101100; b = 8'b11101100; cin = 1'b0; // Expected: {'sum': 152, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101100; b = 8'b11101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1520,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 152, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b10001111; cin = 1'b1; // Expected: {'sum': 139, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b10001111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1521,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 139, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010110; b = 8'b11011001; cin = 1'b1; // Expected: {'sum': 176, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010110; b = 8'b11011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1522,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 176, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000110; b = 8'b11110110; cin = 1'b0; // Expected: {'sum': 188, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000110; b = 8'b11110110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1523,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 188, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b11011110; cin = 1'b0; // Expected: {'sum': 154, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b11011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1524,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 154, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100111; b = 8'b00011010; cin = 1'b0; // Expected: {'sum': 1, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100111; b = 8'b00011010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1525,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b01101100; cin = 1'b1; // Expected: {'sum': 236, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b01101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1526,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 236, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101111; b = 8'b11101010; cin = 1'b1; // Expected: {'sum': 218, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101111; b = 8'b11101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1527,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 218, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b10110011; cin = 1'b1; // Expected: {'sum': 149, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b10110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1528,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 149, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000011; b = 8'b11101010; cin = 1'b1; // Expected: {'sum': 238, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000011; b = 8'b11101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1529,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 238, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b10101011; cin = 1'b0; // Expected: {'sum': 44, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b10101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1530,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 44, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b01011001; cin = 1'b0; // Expected: {'sum': 232, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b01011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1531,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 232, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b01000100; cin = 1'b0; // Expected: {'sum': 252, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b01000100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1532,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 252, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b11010101; cin = 1'b1; // Expected: {'sum': 92, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b11010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1533,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 92, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010100; b = 8'b11110011; cin = 1'b1; // Expected: {'sum': 72, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010100; b = 8'b11110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1534,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 72, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b10101100; cin = 1'b0; // Expected: {'sum': 22, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b10101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1535,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 22, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b01100001; cin = 1'b0; // Expected: {'sum': 73, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b01100001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1536,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 73, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101010; b = 8'b00101110; cin = 1'b1; // Expected: {'sum': 217, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101010; b = 8'b00101110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1537,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 217, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100000; b = 8'b01010000; cin = 1'b1; // Expected: {'sum': 177, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100000; b = 8'b01010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1538,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 177, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b11001101; cin = 1'b1; // Expected: {'sum': 36, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b11001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1539,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 36, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b11100000; cin = 1'b1; // Expected: {'sum': 127, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b11100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1540,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 127, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b10000111; cin = 1'b0; // Expected: {'sum': 37, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b10000111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1541,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 37, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b00000100; cin = 1'b1; // Expected: {'sum': 102, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b00000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1542,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 102, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b10001010; cin = 1'b1; // Expected: {'sum': 118, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b10001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1543,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 118, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b10101101; cin = 1'b1; // Expected: {'sum': 81, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b10101101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1544,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 81, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000011; b = 8'b11100010; cin = 1'b1; // Expected: {'sum': 166, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000011; b = 8'b11100010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1545,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 166, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b11011101; cin = 1'b0; // Expected: {'sum': 74, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b11011101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1546,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 74, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b11011110; cin = 1'b1; // Expected: {'sum': 211, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b11011110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1547,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 211, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001111; b = 8'b10101101; cin = 1'b1; // Expected: {'sum': 189, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001111; b = 8'b10101101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1548,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 189, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010101; b = 8'b10100110; cin = 1'b1; // Expected: {'sum': 188, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010101; b = 8'b10100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1549,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 188, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b01011101; cin = 1'b1; // Expected: {'sum': 70, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b01011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1550,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 70, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b01001001; cin = 1'b1; // Expected: {'sum': 143, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b01001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1551,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 143, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b11111100; cin = 1'b1; // Expected: {'sum': 139, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b11111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1552,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 139, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b01110111; cin = 1'b0; // Expected: {'sum': 104, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b01110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1553,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 104, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b11111010; cin = 1'b0; // Expected: {'sum': 234, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b11111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1554,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 234, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b10100100; cin = 1'b0; // Expected: {'sum': 44, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b10100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1555,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 44, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000100; b = 8'b00101101; cin = 1'b0; // Expected: {'sum': 49, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000100; b = 8'b00101101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1556,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 49, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b01111100; cin = 1'b1; // Expected: {'sum': 97, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b01111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1557,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 97, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b01000100; cin = 1'b0; // Expected: {'sum': 128, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b01000100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1558,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 128, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b10111110; cin = 1'b0; // Expected: {'sum': 99, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b10111110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1559,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 99, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b10000001; cin = 1'b0; // Expected: {'sum': 136, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b10000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1560,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 136, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000011; b = 8'b00001100; cin = 1'b1; // Expected: {'sum': 208, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000011; b = 8'b00001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1561,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 208, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b11110101; cin = 1'b0; // Expected: {'sum': 110, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b11110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1562,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 110, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000101; b = 8'b10010000; cin = 1'b0; // Expected: {'sum': 21, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000101; b = 8'b10010000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1563,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 21, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b11100100; cin = 1'b0; // Expected: {'sum': 98, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b11100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1564,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 98, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b11100000; cin = 1'b0; // Expected: {'sum': 110, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b11100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1565,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 110, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001110; b = 8'b01100011; cin = 1'b0; // Expected: {'sum': 113, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001110; b = 8'b01100011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1566,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 113, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b11110101; cin = 1'b0; // Expected: {'sum': 15, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b11110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1567,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001110; b = 8'b00110110; cin = 1'b1; // Expected: {'sum': 133, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001110; b = 8'b00110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1568,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 133, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101001; b = 8'b01110001; cin = 1'b1; // Expected: {'sum': 91, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101001; b = 8'b01110001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1569,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 91, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b11101111; cin = 1'b0; // Expected: {'sum': 91, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b11101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1570,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 91, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010100; b = 8'b10110000; cin = 1'b0; // Expected: {'sum': 68, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010100; b = 8'b10110000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1571,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 68, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b10010011; cin = 1'b0; // Expected: {'sum': 37, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b10010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1572,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 37, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100000; b = 8'b10100110; cin = 1'b1; // Expected: {'sum': 7, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100000; b = 8'b10100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1573,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b10000110; cin = 1'b1; // Expected: {'sum': 9, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b10000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1574,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 9, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b00011011; cin = 1'b0; // Expected: {'sum': 8, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b00011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1575,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 8, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b01001111; cin = 1'b1; // Expected: {'sum': 79, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b01001111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1576,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 79, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b11100100; cin = 1'b0; // Expected: {'sum': 91, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b11100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1577,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 91, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010100; b = 8'b01000111; cin = 1'b1; // Expected: {'sum': 156, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010100; b = 8'b01000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1578,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 156, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b00001001; cin = 1'b0; // Expected: {'sum': 18, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b00001001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1579,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 18, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b01111010; cin = 1'b1; // Expected: {'sum': 209, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b01111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1580,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 209, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b11110000; cin = 1'b0; // Expected: {'sum': 129, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b11110000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1581,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 129, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100001; b = 8'b00001011; cin = 1'b1; // Expected: {'sum': 45, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100001; b = 8'b00001011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1582,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 45, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000110; b = 8'b10100111; cin = 1'b1; // Expected: {'sum': 238, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000110; b = 8'b10100111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1583,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 238, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b11110100; cin = 1'b0; // Expected: {'sum': 198, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b11110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1584,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 198, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001011; b = 8'b00100011; cin = 1'b1; // Expected: {'sum': 47, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001011; b = 8'b00100011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1585,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 47, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011100; b = 8'b00011000; cin = 1'b0; // Expected: {'sum': 244, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011100; b = 8'b00011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1586,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 244, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b01100010; cin = 1'b0; // Expected: {'sum': 164, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b01100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1587,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 164, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b00001010; cin = 1'b1; // Expected: {'sum': 200, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b00001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1588,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 200, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000110; b = 8'b11010100; cin = 1'b1; // Expected: {'sum': 27, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000110; b = 8'b11010100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1589,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 27, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110101; b = 8'b00000010; cin = 1'b0; // Expected: {'sum': 55, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110101; b = 8'b00000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1590,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 55, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010110; b = 8'b11010010; cin = 1'b0; // Expected: {'sum': 168, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010110; b = 8'b11010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1591,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 168, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010010; b = 8'b11001000; cin = 1'b1; // Expected: {'sum': 27, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010010; b = 8'b11001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1592,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 27, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b11101101; cin = 1'b1; // Expected: {'sum': 148, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b11101101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1593,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 148, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b00011010; cin = 1'b0; // Expected: {'sum': 36, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b00011010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1594,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 36, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000011; b = 8'b00110010; cin = 1'b0; // Expected: {'sum': 245, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000011; b = 8'b00110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1595,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 245, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010011; b = 8'b11011010; cin = 1'b0; // Expected: {'sum': 173, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010011; b = 8'b11011010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1596,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 173, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b10110111; cin = 1'b0; // Expected: {'sum': 250, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b10110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1597,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 250, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b00100100; cin = 1'b0; // Expected: {'sum': 45, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b00100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1598,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 45, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011101; b = 8'b01111101; cin = 1'b1; // Expected: {'sum': 91, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011101; b = 8'b01111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1599,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 91, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b00000100; cin = 1'b1; // Expected: {'sum': 39, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b00000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1600,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 39, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b01011010; cin = 1'b0; // Expected: {'sum': 118, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b01011010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1601,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 118, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101011; b = 8'b00100100; cin = 1'b1; // Expected: {'sum': 80, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101011; b = 8'b00100100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1602,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 80, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b10001000; cin = 1'b0; // Expected: {'sum': 46, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b10001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1603,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 46, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b01001000; cin = 1'b0; // Expected: {'sum': 221, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b01001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1604,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 221, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b11101011; cin = 1'b0; // Expected: {'sum': 167, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b11101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1605,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 167, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001001; b = 8'b01000110; cin = 1'b1; // Expected: {'sum': 144, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001001; b = 8'b01000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1606,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 144, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001101; b = 8'b00000101; cin = 1'b1; // Expected: {'sum': 19, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001101; b = 8'b00000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1607,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 19, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111101; b = 8'b11010100; cin = 1'b0; // Expected: {'sum': 17, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111101; b = 8'b11010100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1608,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 17, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b10111000; cin = 1'b1; // Expected: {'sum': 135, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b10111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1609,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 135, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b01110100; cin = 1'b1; // Expected: {'sum': 168, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b01110100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1610,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 168, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001111; b = 8'b00110111; cin = 1'b0; // Expected: {'sum': 70, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001111; b = 8'b00110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1611,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 70, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b11011101; cin = 1'b0; // Expected: {'sum': 229, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b11011101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1612,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 229, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101111; b = 8'b00000011; cin = 1'b1; // Expected: {'sum': 243, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101111; b = 8'b00000011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1613,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 243, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b01110111; cin = 1'b0; // Expected: {'sum': 32, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b01110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1614,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 32, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b11010100; cin = 1'b0; // Expected: {'sum': 116, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b11010100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1615,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 116, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b10101010; cin = 1'b0; // Expected: {'sum': 198, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b10101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1616,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 198, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001111; b = 8'b01101100; cin = 1'b0; // Expected: {'sum': 187, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001111; b = 8'b01101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1617,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 187, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b11101111; cin = 1'b1; // Expected: {'sum': 94, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b11101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1618,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 94, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110010; b = 8'b11111011; cin = 1'b0; // Expected: {'sum': 109, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110010; b = 8'b11111011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1619,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 109, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b10011001; cin = 1'b0; // Expected: {'sum': 47, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b10011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1620,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 47, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110100; b = 8'b01011000; cin = 1'b1; // Expected: {'sum': 205, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110100; b = 8'b01011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1621,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 205, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b11011000; cin = 1'b1; // Expected: {'sum': 106, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b11011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1622,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 106, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b11101010; cin = 1'b1; // Expected: {'sum': 185, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b11101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1623,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 185, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b00001011; cin = 1'b1; // Expected: {'sum': 142, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b00001011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1624,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 142, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b01111001; cin = 1'b0; // Expected: {'sum': 252, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b01111001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1625,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 252, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b00100010; cin = 1'b1; // Expected: {'sum': 58, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b00100010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1626,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 58, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111001; b = 8'b01100000; cin = 1'b0; // Expected: {'sum': 153, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111001; b = 8'b01100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1627,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 153, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100010; b = 8'b11011110; cin = 1'b0; // Expected: {'sum': 128, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100010; b = 8'b11011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1628,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 128, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b01000101; cin = 1'b1; // Expected: {'sum': 43, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b01000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1629,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 43, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000011; b = 8'b11011111; cin = 1'b0; // Expected: {'sum': 226, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000011; b = 8'b11011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1630,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 226, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b11101100; cin = 1'b1; // Expected: {'sum': 31, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b11101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1631,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 31, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100000; b = 8'b01010100; cin = 1'b0; // Expected: {'sum': 52, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100000; b = 8'b01010100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1632,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 52, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100111; b = 8'b00111101; cin = 1'b1; // Expected: {'sum': 229, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100111; b = 8'b00111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1633,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 229, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b00110101; cin = 1'b1; // Expected: {'sum': 21, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b00110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1634,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 21, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b11101001; cin = 1'b1; // Expected: {'sum': 87, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b11101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1635,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 87, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b11011010; cin = 1'b1; // Expected: {'sum': 27, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b11011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1636,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 27, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000111; b = 8'b01100001; cin = 1'b0; // Expected: {'sum': 232, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000111; b = 8'b01100001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1637,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 232, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b00101010; cin = 1'b1; // Expected: {'sum': 211, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b00101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1638,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 211, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b01011001; cin = 1'b0; // Expected: {'sum': 112, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b01011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1639,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 112, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b10110100; cin = 1'b0; // Expected: {'sum': 130, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b10110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1640,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 130, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001100; b = 8'b11101101; cin = 1'b0; // Expected: {'sum': 249, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001100; b = 8'b11101101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1641,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 249, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b11010110; cin = 1'b0; // Expected: {'sum': 193, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b11010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1642,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 193, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b10111100; cin = 1'b0; // Expected: {'sum': 3, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b10111100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1643,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011101; b = 8'b00110010; cin = 1'b0; // Expected: {'sum': 15, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011101; b = 8'b00110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1644,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101110; b = 8'b01011010; cin = 1'b0; // Expected: {'sum': 8, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101110; b = 8'b01011010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1645,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 8, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000011; b = 8'b01100100; cin = 1'b1; // Expected: {'sum': 40, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000011; b = 8'b01100100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1646,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 40, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b01000111; cin = 1'b1; // Expected: {'sum': 58, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b01000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1647,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 58, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011011; b = 8'b10110100; cin = 1'b1; // Expected: {'sum': 208, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011011; b = 8'b10110100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1648,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 208, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b11111101; cin = 1'b0; // Expected: {'sum': 7, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b11111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1649,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b10000111; cin = 1'b0; // Expected: {'sum': 215, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b10000111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1650,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 215, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000011; b = 8'b10111001; cin = 1'b1; // Expected: {'sum': 125, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000011; b = 8'b10111001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1651,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 125, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b11011111; cin = 1'b0; // Expected: {'sum': 232, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b11011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1652,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 232, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100010; b = 8'b00111101; cin = 1'b1; // Expected: {'sum': 32, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100010; b = 8'b00111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1653,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 32, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b10101000; cin = 1'b1; // Expected: {'sum': 123, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b10101000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1654,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 123, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b00001011; cin = 1'b0; // Expected: {'sum': 224, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b00001011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1655,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 224, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011101; b = 8'b00010011; cin = 1'b1; // Expected: {'sum': 241, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011101; b = 8'b00010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1656,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 241, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b00100011; cin = 1'b0; // Expected: {'sum': 87, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b00100011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1657,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 87, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b11001011; cin = 1'b1; // Expected: {'sum': 54, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b11001011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1658,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 54, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b00001001; cin = 1'b0; // Expected: {'sum': 129, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b00001001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1659,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 129, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b01010011; cin = 1'b1; // Expected: {'sum': 225, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b01010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1660,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 225, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000110; b = 8'b10010000; cin = 1'b1; // Expected: {'sum': 215, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000110; b = 8'b10010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1661,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 215, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b11000010; cin = 1'b1; // Expected: {'sum': 158, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b11000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1662,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 158, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110000; b = 8'b10111000; cin = 1'b1; // Expected: {'sum': 233, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110000; b = 8'b10111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1663,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 233, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111000; b = 8'b00010100; cin = 1'b0; // Expected: {'sum': 12, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111000; b = 8'b00010100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1664,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b00101100; cin = 1'b0; // Expected: {'sum': 79, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b00101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1665,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 79, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001100; b = 8'b00010101; cin = 1'b0; // Expected: {'sum': 161, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001100; b = 8'b00010101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1666,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 161, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b01110000; cin = 1'b0; // Expected: {'sum': 63, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b01110000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1667,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 63, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100000; b = 8'b00111010; cin = 1'b1; // Expected: {'sum': 91, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100000; b = 8'b00111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1668,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 91, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b00000001; cin = 1'b1; // Expected: {'sum': 66, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b00000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1669,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 66, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000101; b = 8'b10001101; cin = 1'b1; // Expected: {'sum': 19, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000101; b = 8'b10001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1670,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 19, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b10000011; cin = 1'b1; // Expected: {'sum': 156, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b10000011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1671,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 156, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110110; b = 8'b00010110; cin = 1'b0; // Expected: {'sum': 140, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110110; b = 8'b00010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1672,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 140, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100110; b = 8'b10110001; cin = 1'b0; // Expected: {'sum': 215, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100110; b = 8'b10110001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1673,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 215, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010111; b = 8'b00010001; cin = 1'b0; // Expected: {'sum': 104, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010111; b = 8'b00010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1674,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 104, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b11000110; cin = 1'b0; // Expected: {'sum': 227, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b11000110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1675,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 227, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b10111010; cin = 1'b1; // Expected: {'sum': 74, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b10111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1676,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 74, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110100; b = 8'b11101111; cin = 1'b1; // Expected: {'sum': 100, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110100; b = 8'b11101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1677,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 100, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b11101101; cin = 1'b0; // Expected: {'sum': 139, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b11101101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1678,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 139, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b10010101; cin = 1'b1; // Expected: {'sum': 158, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b10010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1679,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 158, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001111; b = 8'b10010000; cin = 1'b0; // Expected: {'sum': 223, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001111; b = 8'b10010000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1680,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 223, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b11001011; cin = 1'b1; // Expected: {'sum': 221, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b11001011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1681,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 221, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b11001010; cin = 1'b0; // Expected: {'sum': 197, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b11001010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1682,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 197, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b00001100; cin = 1'b0; // Expected: {'sum': 57, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b00001100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1683,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 57, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010100; b = 8'b01100000; cin = 1'b0; // Expected: {'sum': 244, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010100; b = 8'b01100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1684,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 244, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b01100100; cin = 1'b1; // Expected: {'sum': 52, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b01100100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1685,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 52, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101010; b = 8'b01101011; cin = 1'b1; // Expected: {'sum': 86, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101010; b = 8'b01101011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1686,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 86, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b00110010; cin = 1'b1; // Expected: {'sum': 227, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b00110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1687,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 227, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b00100010; cin = 1'b1; // Expected: {'sum': 112, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b00100010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1688,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 112, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b00101111; cin = 1'b0; // Expected: {'sum': 249, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b00101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1689,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 249, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b00001101; cin = 1'b0; // Expected: {'sum': 80, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b00001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1690,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 80, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100001; b = 8'b00001100; cin = 1'b1; // Expected: {'sum': 46, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100001; b = 8'b00001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1691,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 46, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b01011110; cin = 1'b0; // Expected: {'sum': 94, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b01011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1692,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 94, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011010; b = 8'b01011111; cin = 1'b1; // Expected: {'sum': 250, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011010; b = 8'b01011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1693,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 250, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b10010100; cin = 1'b0; // Expected: {'sum': 50, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b10010100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1694,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 50, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001011; b = 8'b10101011; cin = 1'b1; // Expected: {'sum': 247, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001011; b = 8'b10101011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1695,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 247, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b10010011; cin = 1'b0; // Expected: {'sum': 49, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b10010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1696,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 49, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b11000101; cin = 1'b1; // Expected: {'sum': 128, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b11000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1697,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 128, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010100; b = 8'b10110100; cin = 1'b0; // Expected: {'sum': 136, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010100; b = 8'b10110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1698,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 136, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b10010100; cin = 1'b1; // Expected: {'sum': 128, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b10010100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1699,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 128, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101111; b = 8'b11111111; cin = 1'b1; // Expected: {'sum': 239, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101111; b = 8'b11111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1700,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 239, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b01000010; cin = 1'b1; // Expected: {'sum': 218, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b01000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1701,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 218, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b11101110; cin = 1'b0; // Expected: {'sum': 36, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b11101110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1702,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 36, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b11101011; cin = 1'b1; // Expected: {'sum': 199, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b11101011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1703,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 199, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100111; b = 8'b11101100; cin = 1'b1; // Expected: {'sum': 212, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100111; b = 8'b11101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1704,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 212, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010010; b = 8'b01110010; cin = 1'b0; // Expected: {'sum': 196, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010010; b = 8'b01110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1705,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 196, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b11001100; cin = 1'b1; // Expected: {'sum': 57, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b11001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1706,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 57, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b10100110; cin = 1'b1; // Expected: {'sum': 244, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b10100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1707,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 244, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b01101100; cin = 1'b1; // Expected: {'sum': 95, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b01101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1708,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 95, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001011; b = 8'b10101110; cin = 1'b1; // Expected: {'sum': 122, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001011; b = 8'b10101110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1709,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 122, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100001; b = 8'b11010111; cin = 1'b1; // Expected: {'sum': 249, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100001; b = 8'b11010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1710,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 249, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b00001101; cin = 1'b1; // Expected: {'sum': 95, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b00001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1711,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 95, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b01111101; cin = 1'b0; // Expected: {'sum': 226, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b01111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1712,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 226, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001111; b = 8'b11100111; cin = 1'b1; // Expected: {'sum': 55, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001111; b = 8'b11100111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1713,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 55, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010010; b = 8'b10001110; cin = 1'b1; // Expected: {'sum': 225, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010010; b = 8'b10001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1714,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 225, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110000; b = 8'b01100010; cin = 1'b1; // Expected: {'sum': 147, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110000; b = 8'b01100010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1715,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 147, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000111; b = 8'b01100010; cin = 1'b1; // Expected: {'sum': 234, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000111; b = 8'b01100010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1716,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 234, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b10011001; cin = 1'b1; // Expected: {'sum': 106, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b10011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1717,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 106, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b10100100; cin = 1'b1; // Expected: {'sum': 58, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b10100100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1718,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 58, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b11001000; cin = 1'b0; // Expected: {'sum': 95, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b11001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1719,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 95, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b00100010; cin = 1'b0; // Expected: {'sum': 44, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b00100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1720,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 44, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b11110001; cin = 1'b0; // Expected: {'sum': 193, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b11110001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1721,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 193, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101010; b = 8'b11111010; cin = 1'b1; // Expected: {'sum': 165, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101010; b = 8'b11111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1722,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 165, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b01110000; cin = 1'b1; // Expected: {'sum': 250, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b01110000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1723,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 250, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b10000010; cin = 1'b0; // Expected: {'sum': 216, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b10000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1724,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 216, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b00010010; cin = 1'b1; // Expected: {'sum': 123, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b00010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1725,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 123, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010101; b = 8'b01110011; cin = 1'b1; // Expected: {'sum': 137, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010101; b = 8'b01110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1726,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 137, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000011; b = 8'b11011010; cin = 1'b1; // Expected: {'sum': 158, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000011; b = 8'b11011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1727,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 158, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b10010101; cin = 1'b0; // Expected: {'sum': 118, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b10010101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1728,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 118, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010101; b = 8'b01010000; cin = 1'b1; // Expected: {'sum': 102, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010101; b = 8'b01010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1729,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 102, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110010; b = 8'b10110010; cin = 1'b1; // Expected: {'sum': 37, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110010; b = 8'b10110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1730,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 37, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b00100000; cin = 1'b0; // Expected: {'sum': 25, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b00100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1731,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 25, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b10011101; cin = 1'b0; // Expected: {'sum': 129, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b10011101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1732,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 129, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100010; b = 8'b01101001; cin = 1'b0; // Expected: {'sum': 75, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100010; b = 8'b01101001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1733,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 75, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b00101001; cin = 1'b0; // Expected: {'sum': 233, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b00101001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1734,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 233, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b10100110; cin = 1'b1; // Expected: {'sum': 105, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b10100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1735,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 105, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b00010101; cin = 1'b1; // Expected: {'sum': 143, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b00010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1736,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 143, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b01001010; cin = 1'b0; // Expected: {'sum': 154, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b01001010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1737,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 154, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b11001110; cin = 1'b1; // Expected: {'sum': 28, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b11001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1738,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 28, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b00010011; cin = 1'b0; // Expected: {'sum': 28, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b00010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1739,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 28, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b01111000; cin = 1'b0; // Expected: {'sum': 241, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b01111000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1740,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 241, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101111; b = 8'b01101000; cin = 1'b0; // Expected: {'sum': 87, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101111; b = 8'b01101000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1741,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 87, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b01100111; cin = 1'b0; // Expected: {'sum': 132, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b01100111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1742,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 132, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b00000001; cin = 1'b0; // Expected: {'sum': 128, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b00000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1743,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 128, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b10100111; cin = 1'b1; // Expected: {'sum': 61, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b10100111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1744,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 61, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101001; b = 8'b10101010; cin = 1'b1; // Expected: {'sum': 20, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101001; b = 8'b10101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1745,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 20, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b01110011; cin = 1'b1; // Expected: {'sum': 54, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b01110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1746,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 54, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b11011011; cin = 1'b0; // Expected: {'sum': 109, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b11011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1747,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 109, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011100; b = 8'b00000101; cin = 1'b1; // Expected: {'sum': 226, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011100; b = 8'b00000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1748,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 226, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010100; b = 8'b10111000; cin = 1'b1; // Expected: {'sum': 141, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010100; b = 8'b10111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1749,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 141, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010001; b = 8'b11001011; cin = 1'b1; // Expected: {'sum': 157, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010001; b = 8'b11001011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1750,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 157, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100010; b = 8'b10011011; cin = 1'b1; // Expected: {'sum': 62, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100010; b = 8'b10011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1751,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 62, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101111; b = 8'b01100001; cin = 1'b1; // Expected: {'sum': 209, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101111; b = 8'b01100001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1752,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 209, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011010; b = 8'b01100101; cin = 1'b0; // Expected: {'sum': 191, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011010; b = 8'b01100101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1753,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 191, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b00111010; cin = 1'b1; // Expected: {'sum': 111, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b00111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1754,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 111, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b10001011; cin = 1'b1; // Expected: {'sum': 237, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b10001011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1755,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 237, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b00001101; cin = 1'b0; // Expected: {'sum': 202, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b00001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1756,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 202, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b00001111; cin = 1'b1; // Expected: {'sum': 117, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b00001111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1757,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 117, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010100; b = 8'b01110001; cin = 1'b1; // Expected: {'sum': 198, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010100; b = 8'b01110001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1758,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 198, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100001; b = 8'b10111000; cin = 1'b1; // Expected: {'sum': 218, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100001; b = 8'b10111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1759,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 218, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001110; b = 8'b01110011; cin = 1'b1; // Expected: {'sum': 194, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001110; b = 8'b01110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1760,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 194, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b00001011; cin = 1'b1; // Expected: {'sum': 156, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b00001011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1761,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 156, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100010; b = 8'b00011110; cin = 1'b0; // Expected: {'sum': 192, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100010; b = 8'b00011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1762,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 192, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b11011001; cin = 1'b1; // Expected: {'sum': 148, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b11011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1763,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 148, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b11111101; cin = 1'b0; // Expected: {'sum': 234, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b11111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1764,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 234, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101111; b = 8'b00001011; cin = 1'b1; // Expected: {'sum': 251, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101111; b = 8'b00001011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1765,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 251, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b00010110; cin = 1'b1; // Expected: {'sum': 31, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b00010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1766,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 31, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b00000010; cin = 1'b1; // Expected: {'sum': 80, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b00000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1767,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 80, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b01010010; cin = 1'b1; // Expected: {'sum': 152, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b01010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1768,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 152, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b00110011; cin = 1'b0; // Expected: {'sum': 144, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b00110011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1769,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 144, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011000; b = 8'b10010011; cin = 1'b1; // Expected: {'sum': 236, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011000; b = 8'b10010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1770,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 236, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b00010010; cin = 1'b0; // Expected: {'sum': 133, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b00010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1771,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 133, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101110; b = 8'b10110011; cin = 1'b1; // Expected: {'sum': 98, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101110; b = 8'b10110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1772,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 98, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110001; b = 8'b00000111; cin = 1'b1; // Expected: {'sum': 121, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110001; b = 8'b00000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1773,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 121, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011010; b = 8'b00011010; cin = 1'b0; // Expected: {'sum': 244, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011010; b = 8'b00011010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1774,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 244, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001110; b = 8'b01011011; cin = 1'b1; // Expected: {'sum': 170, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001110; b = 8'b01011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1775,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 170, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b00111011; cin = 1'b0; // Expected: {'sum': 202, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b00111011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1776,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 202, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b10110110; cin = 1'b0; // Expected: {'sum': 206, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b10110110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1777,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 206, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b11111000; cin = 1'b0; // Expected: {'sum': 96, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b11111000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1778,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 96, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b01100101; cin = 1'b1; // Expected: {'sum': 84, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b01100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1779,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 84, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010011; b = 8'b10000010; cin = 1'b0; // Expected: {'sum': 85, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010011; b = 8'b10000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1780,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 85, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b10011000; cin = 1'b1; // Expected: {'sum': 52, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b10011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1781,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 52, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b00101100; cin = 1'b0; // Expected: {'sum': 148, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b00101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1782,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 148, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b01101010; cin = 1'b1; // Expected: {'sum': 66, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b01101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1783,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 66, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b10010101; cin = 1'b1; // Expected: {'sum': 227, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b10010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1784,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 227, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101101; b = 8'b00111111; cin = 1'b1; // Expected: {'sum': 237, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101101; b = 8'b00111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1785,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 237, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b00000001; cin = 1'b1; // Expected: {'sum': 204, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b00000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1786,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 204, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b01100011; cin = 1'b0; // Expected: {'sum': 51, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b01100011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1787,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 51, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b10011101; cin = 1'b1; // Expected: {'sum': 62, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b10011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1788,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 62, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111011; b = 8'b11111011; cin = 1'b1; // Expected: {'sum': 119, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111011; b = 8'b11111011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1789,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 119, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101100; b = 8'b00110101; cin = 1'b1; // Expected: {'sum': 34, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101100; b = 8'b00110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1790,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 34, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100110; b = 8'b00011010; cin = 1'b1; // Expected: {'sum': 129, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100110; b = 8'b00011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1791,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 129, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101010; b = 8'b10000001; cin = 1'b0; // Expected: {'sum': 171, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101010; b = 8'b10000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1792,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 171, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111000; b = 8'b10011111; cin = 1'b0; // Expected: {'sum': 151, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111000; b = 8'b10011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1793,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 151, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b10110001; cin = 1'b0; // Expected: {'sum': 170, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b10110001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1794,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 170, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b00111100; cin = 1'b0; // Expected: {'sum': 210, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b00111100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1795,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 210, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b01010110; cin = 1'b0; // Expected: {'sum': 236, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b01010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1796,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 236, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b00110010; cin = 1'b0; // Expected: {'sum': 4, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b00110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1797,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001101; b = 8'b10101111; cin = 1'b1; // Expected: {'sum': 189, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001101; b = 8'b10101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1798,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 189, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b01011001; cin = 1'b0; // Expected: {'sum': 196, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b01011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1799,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 196, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b01010111; cin = 1'b0; // Expected: {'sum': 88, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b01010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1800,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 88, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b01111100; cin = 1'b1; // Expected: {'sum': 14, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b01111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1801,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b11111101; cin = 1'b1; // Expected: {'sum': 69, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b11111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1802,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 69, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110110; b = 8'b01011001; cin = 1'b0; // Expected: {'sum': 207, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110110; b = 8'b01011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1803,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 207, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b00111101; cin = 1'b0; // Expected: {'sum': 217, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b00111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1804,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 217, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011110; b = 8'b11000100; cin = 1'b1; // Expected: {'sum': 163, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011110; b = 8'b11000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1805,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 163, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101111; b = 8'b01010110; cin = 1'b1; // Expected: {'sum': 198, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101111; b = 8'b01010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1806,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 198, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b10011011; cin = 1'b0; // Expected: {'sum': 35, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b10011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1807,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 35, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101010; b = 8'b00111010; cin = 1'b0; // Expected: {'sum': 36, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101010; b = 8'b00111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1808,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 36, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b00001100; cin = 1'b0; // Expected: {'sum': 70, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b00001100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1809,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 70, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b01111000; cin = 1'b1; // Expected: {'sum': 188, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b01111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1810,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 188, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101100; b = 8'b00000100; cin = 1'b0; // Expected: {'sum': 176, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101100; b = 8'b00000100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1811,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 176, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b01010111; cin = 1'b1; // Expected: {'sum': 88, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b01010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1812,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 88, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b10001110; cin = 1'b1; // Expected: {'sum': 212, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b10001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1813,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 212, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b01001011; cin = 1'b1; // Expected: {'sum': 39, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b01001011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1814,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 39, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b00101100; cin = 1'b0; // Expected: {'sum': 96, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b00101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1815,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 96, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b11001111; cin = 1'b0; // Expected: {'sum': 11, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b11001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1816,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 11, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b10100010; cin = 1'b0; // Expected: {'sum': 125, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b10100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1817,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 125, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b10101110; cin = 1'b0; // Expected: {'sum': 60, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b10101110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1818,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 60, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b11010110; cin = 1'b0; // Expected: {'sum': 249, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b11010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1819,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 249, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b00000011; cin = 1'b1; // Expected: {'sum': 146, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b00000011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1820,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 146, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b10110101; cin = 1'b0; // Expected: {'sum': 55, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b10110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1821,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 55, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010100; b = 8'b01111100; cin = 1'b0; // Expected: {'sum': 80, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010100; b = 8'b01111100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1822,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 80, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b01100110; cin = 1'b0; // Expected: {'sum': 130, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b01100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1823,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 130, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b10001100; cin = 1'b0; // Expected: {'sum': 10, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b10001100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1824,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b01001000; cin = 1'b0; // Expected: {'sum': 176, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b01001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1825,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 176, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b00100100; cin = 1'b0; // Expected: {'sum': 27, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b00100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1826,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 27, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001111; b = 8'b10101011; cin = 1'b0; // Expected: {'sum': 250, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001111; b = 8'b10101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1827,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 250, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b00001110; cin = 1'b1; // Expected: {'sum': 146, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b00001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1828,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 146, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b01010001; cin = 1'b0; // Expected: {'sum': 217, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b01010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1829,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 217, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100001; b = 8'b00111110; cin = 1'b0; // Expected: {'sum': 95, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100001; b = 8'b00111110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1830,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 95, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b10010101; cin = 1'b0; // Expected: {'sum': 82, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b10010101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1831,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 82, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001111; b = 8'b01111000; cin = 1'b1; // Expected: {'sum': 200, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001111; b = 8'b01111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1832,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 200, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111101; b = 8'b00110110; cin = 1'b1; // Expected: {'sum': 52, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111101; b = 8'b00110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1833,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 52, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b01010101; cin = 1'b1; // Expected: {'sum': 120, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b01010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1834,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 120, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b01001110; cin = 1'b1; // Expected: {'sum': 51, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b01001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1835,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 51, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b10110110; cin = 1'b1; // Expected: {'sum': 137, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b10110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1836,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 137, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111000; b = 8'b00010000; cin = 1'b0; // Expected: {'sum': 72, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111000; b = 8'b00010000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1837,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 72, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010011; b = 8'b01111010; cin = 1'b1; // Expected: {'sum': 206, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010011; b = 8'b01111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1838,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 206, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b00111101; cin = 1'b0; // Expected: {'sum': 57, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b00111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1839,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 57, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b01100010; cin = 1'b1; // Expected: {'sum': 245, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b01100010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1840,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 245, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b10101010; cin = 1'b0; // Expected: {'sum': 85, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b10101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1841,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 85, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b01110100; cin = 1'b0; // Expected: {'sum': 45, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b01110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1842,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 45, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100111; b = 8'b00101001; cin = 1'b1; // Expected: {'sum': 145, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100111; b = 8'b00101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1843,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 145, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111111; b = 8'b11010110; cin = 1'b0; // Expected: {'sum': 21, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111111; b = 8'b11010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1844,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 21, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b11100001; cin = 1'b1; // Expected: {'sum': 128, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b11100001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1845,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 128, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b11011110; cin = 1'b0; // Expected: {'sum': 121, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b11011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1846,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 121, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010100; b = 8'b01000111; cin = 1'b1; // Expected: {'sum': 28, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010100; b = 8'b01000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1847,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 28, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b01101001; cin = 1'b1; // Expected: {'sum': 248, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b01101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1848,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 248, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110000; b = 8'b10010010; cin = 1'b1; // Expected: {'sum': 3, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110000; b = 8'b10010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1849,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b00001000; cin = 1'b1; // Expected: {'sum': 216, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b00001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1850,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 216, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b00000011; cin = 1'b1; // Expected: {'sum': 217, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b00000011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1851,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 217, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110000; b = 8'b01000000; cin = 1'b0; // Expected: {'sum': 112, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110000; b = 8'b01000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1852,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 112, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010011; b = 8'b10001000; cin = 1'b1; // Expected: {'sum': 92, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010011; b = 8'b10001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1853,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 92, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b10110110; cin = 1'b0; // Expected: {'sum': 36, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b10110110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1854,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 36, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b00101101; cin = 1'b0; // Expected: {'sum': 153, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b00101101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1855,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 153, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b10110111; cin = 1'b1; // Expected: {'sum': 22, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b10110111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1856,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 22, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010101; b = 8'b11101110; cin = 1'b1; // Expected: {'sum': 68, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010101; b = 8'b11101110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1857,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 68, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000100; b = 8'b01111101; cin = 1'b0; // Expected: {'sum': 129, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000100; b = 8'b01111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1858,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 129, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b01101001; cin = 1'b1; // Expected: {'sum': 111, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b01101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1859,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 111, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b11101000; cin = 1'b1; // Expected: {'sum': 161, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b11101000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1860,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 161, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000101; b = 8'b00010000; cin = 1'b0; // Expected: {'sum': 149, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000101; b = 8'b00010000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1861,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 149, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b11111011; cin = 1'b1; // Expected: {'sum': 239, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b11111011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1862,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 239, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000110; b = 8'b11110001; cin = 1'b0; // Expected: {'sum': 247, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000110; b = 8'b11110001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1863,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 247, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011111; b = 8'b01101110; cin = 1'b0; // Expected: {'sum': 13, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011111; b = 8'b01101110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1864,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 13, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101100; b = 8'b10001001; cin = 1'b1; // Expected: {'sum': 118, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101100; b = 8'b10001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1865,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 118, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b11001111; cin = 1'b0; // Expected: {'sum': 131, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b11001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1866,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 131, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b01010011; cin = 1'b0; // Expected: {'sum': 239, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b01010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1867,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 239, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b01110010; cin = 1'b1; // Expected: {'sum': 78, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b01110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1868,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 78, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b11111001; cin = 1'b1; // Expected: {'sum': 128, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b11111001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1869,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 128, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b10110101; cin = 1'b0; // Expected: {'sum': 176, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b10110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1870,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 176, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b10111111; cin = 1'b1; // Expected: {'sum': 149, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b10111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1871,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 149, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b00011110; cin = 1'b1; // Expected: {'sum': 248, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b00011110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1872,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 248, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b01111011; cin = 1'b1; // Expected: {'sum': 44, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b01111011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1873,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 44, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b10001010; cin = 1'b1; // Expected: {'sum': 233, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b10001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1874,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 233, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b11011011; cin = 1'b0; // Expected: {'sum': 198, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b11011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1875,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 198, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b10110010; cin = 1'b1; // Expected: {'sum': 31, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b10110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1876,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 31, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b00001010; cin = 1'b0; // Expected: {'sum': 173, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b00001010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1877,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 173, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b00100011; cin = 1'b1; // Expected: {'sum': 226, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b00100011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1878,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 226, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b11011010; cin = 1'b1; // Expected: {'sum': 178, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b11011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1879,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 178, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b01110010; cin = 1'b1; // Expected: {'sum': 0, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b01110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1880,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b00101010; cin = 1'b0; // Expected: {'sum': 140, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b00101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1881,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 140, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110101; b = 8'b11011011; cin = 1'b1; // Expected: {'sum': 145, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110101; b = 8'b11011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1882,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 145, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b01000110; cin = 1'b1; // Expected: {'sum': 66, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b01000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1883,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 66, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101001; b = 8'b10100110; cin = 1'b1; // Expected: {'sum': 144, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101001; b = 8'b10100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1884,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 144, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b01101100; cin = 1'b0; // Expected: {'sum': 125, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b01101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1885,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 125, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b01000111; cin = 1'b1; // Expected: {'sum': 139, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b01000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1886,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 139, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b01000110; cin = 1'b1; // Expected: {'sum': 254, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b01000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1887,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 254, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b01010011; cin = 1'b0; // Expected: {'sum': 182, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b01010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1888,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 182, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101111; b = 8'b10100101; cin = 1'b1; // Expected: {'sum': 149, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101111; b = 8'b10100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1889,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 149, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b01110101; cin = 1'b1; // Expected: {'sum': 68, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b01110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1890,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 68, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b00010110; cin = 1'b1; // Expected: {'sum': 148, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b00010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1891,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 148, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b00000010; cin = 1'b1; // Expected: {'sum': 209, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b00000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1892,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 209, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010111; b = 8'b10101100; cin = 1'b1; // Expected: {'sum': 4, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010111; b = 8'b10101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1893,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b01111010; cin = 1'b0; // Expected: {'sum': 55, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b01111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1894,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 55, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b00110010; cin = 1'b1; // Expected: {'sum': 46, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b00110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1895,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 46, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110010; b = 8'b01111010; cin = 1'b0; // Expected: {'sum': 236, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110010; b = 8'b01111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1896,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 236, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011111; b = 8'b11001010; cin = 1'b0; // Expected: {'sum': 41, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011111; b = 8'b11001010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1897,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 41, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b01010000; cin = 1'b0; // Expected: {'sum': 9, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b01010000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1898,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 9, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101100; b = 8'b10000001; cin = 1'b1; // Expected: {'sum': 46, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101100; b = 8'b10000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1899,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 46, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100110; b = 8'b11010011; cin = 1'b0; // Expected: {'sum': 57, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100110; b = 8'b11010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1900,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 57, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010011; b = 8'b01101001; cin = 1'b0; // Expected: {'sum': 252, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010011; b = 8'b01101001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1901,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 252, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b11110100; cin = 1'b0; // Expected: {'sum': 97, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b11110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1902,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 97, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b01101111; cin = 1'b0; // Expected: {'sum': 21, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b01101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1903,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 21, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b00110010; cin = 1'b0; // Expected: {'sum': 35, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b00110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1904,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 35, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010111; b = 8'b01001011; cin = 1'b1; // Expected: {'sum': 163, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010111; b = 8'b01001011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1905,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 163, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b01100100; cin = 1'b1; // Expected: {'sum': 146, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b01100100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1906,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 146, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110110; b = 8'b10111011; cin = 1'b1; // Expected: {'sum': 50, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110110; b = 8'b10111011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1907,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 50, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000111; b = 8'b00100000; cin = 1'b0; // Expected: {'sum': 231, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000111; b = 8'b00100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1908,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 231, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101010; b = 8'b11001010; cin = 1'b1; // Expected: {'sum': 245, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101010; b = 8'b11001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1909,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 245, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b10111111; cin = 1'b1; // Expected: {'sum': 94, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b10111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1910,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 94, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b10001001; cin = 1'b1; // Expected: {'sum': 60, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b10001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1911,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 60, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b11010110; cin = 1'b1; // Expected: {'sum': 59, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b11010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1912,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 59, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b10100011; cin = 1'b1; // Expected: {'sum': 42, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b10100011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1913,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 42, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b11011101; cin = 1'b0; // Expected: {'sum': 208, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b11011101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1914,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 208, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b11101110; cin = 1'b0; // Expected: {'sum': 123, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b11101110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1915,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 123, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b00101011; cin = 1'b0; // Expected: {'sum': 211, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b00101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1916,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 211, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100100; b = 8'b00011110; cin = 1'b0; // Expected: {'sum': 194, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100100; b = 8'b00011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1917,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 194, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b01001100; cin = 1'b1; // Expected: {'sum': 127, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b01001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1918,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 127, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b00000010; cin = 1'b1; // Expected: {'sum': 31, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b00000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1919,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 31, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011001; b = 8'b00000100; cin = 1'b1; // Expected: {'sum': 158, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011001; b = 8'b00000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1920,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 158, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b10110110; cin = 1'b1; // Expected: {'sum': 200, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b10110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1921,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 200, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b11101010; cin = 1'b1; // Expected: {'sum': 56, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b11101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1922,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 56, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011110; b = 8'b00001110; cin = 1'b1; // Expected: {'sum': 237, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011110; b = 8'b00001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1923,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 237, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b00101000; cin = 1'b1; // Expected: {'sum': 78, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b00101000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1924,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 78, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001110; b = 8'b11001000; cin = 1'b0; // Expected: {'sum': 22, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001110; b = 8'b11001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1925,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 22, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b01100001; cin = 1'b1; // Expected: {'sum': 99, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b01100001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1926,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 99, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b01000011; cin = 1'b0; // Expected: {'sum': 49, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b01000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1927,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 49, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110110; b = 8'b11001011; cin = 1'b1; // Expected: {'sum': 66, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110110; b = 8'b11001011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1928,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 66, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b00101011; cin = 1'b1; // Expected: {'sum': 170, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b00101011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1929,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 170, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101011; b = 8'b01010010; cin = 1'b0; // Expected: {'sum': 125, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101011; b = 8'b01010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1930,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 125, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b01000110; cin = 1'b1; // Expected: {'sum': 64, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b01000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1931,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 64, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011001; b = 8'b10100011; cin = 1'b0; // Expected: {'sum': 188, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011001; b = 8'b10100011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1932,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 188, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b01001101; cin = 1'b0; // Expected: {'sum': 7, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b01001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1933,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100000; b = 8'b10110000; cin = 1'b0; // Expected: {'sum': 208, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100000; b = 8'b10110000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1934,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 208, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b00101111; cin = 1'b0; // Expected: {'sum': 101, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b00101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1935,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 101, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b01101110; cin = 1'b1; // Expected: {'sum': 113, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b01101110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1936,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 113, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010101; b = 8'b10011011; cin = 1'b0; // Expected: {'sum': 240, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010101; b = 8'b10011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1937,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 240, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b01110111; cin = 1'b0; // Expected: {'sum': 24, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b01110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1938,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 24, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b00011001; cin = 1'b1; // Expected: {'sum': 106, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b00011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1939,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 106, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b00001111; cin = 1'b1; // Expected: {'sum': 4, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b00001111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1940,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b11110011; cin = 1'b1; // Expected: {'sum': 12, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b11110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1941,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110001; b = 8'b00000111; cin = 1'b1; // Expected: {'sum': 57, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110001; b = 8'b00000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1942,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 57, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b11100111; cin = 1'b1; // Expected: {'sum': 231, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b11100111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1943,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 231, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010101; b = 8'b00101111; cin = 1'b1; // Expected: {'sum': 69, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010101; b = 8'b00101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1944,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 69, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000001; b = 8'b10001000; cin = 1'b1; // Expected: {'sum': 74, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000001; b = 8'b10001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1945,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 74, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b11100100; cin = 1'b1; // Expected: {'sum': 159, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b11100100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1946,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 159, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b01100010; cin = 1'b1; // Expected: {'sum': 216, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b01100010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1947,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 216, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b11100001; cin = 1'b1; // Expected: {'sum': 111, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b11100001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1948,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 111, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b11010001; cin = 1'b0; // Expected: {'sum': 136, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b11010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1949,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 136, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b10001111; cin = 1'b0; // Expected: {'sum': 150, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b10001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1950,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 150, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000110; b = 8'b01111010; cin = 1'b0; // Expected: {'sum': 128, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000110; b = 8'b01111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1951,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 128, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b00000100; cin = 1'b1; // Expected: {'sum': 222, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b00000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1952,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 222, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b10011101; cin = 1'b1; // Expected: {'sum': 71, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b10011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1953,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 71, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b01100101; cin = 1'b1; // Expected: {'sum': 26, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b01100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1954,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 26, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010110; b = 8'b11101010; cin = 1'b1; // Expected: {'sum': 193, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010110; b = 8'b11101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1955,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 193, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b10011011; cin = 1'b1; // Expected: {'sum': 31, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b10011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1956,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 31, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111000; b = 8'b01010000; cin = 1'b0; // Expected: {'sum': 72, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111000; b = 8'b01010000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1957,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 72, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111011; b = 8'b11111000; cin = 1'b0; // Expected: {'sum': 51, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111011; b = 8'b11111000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1958,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 51, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b10001111; cin = 1'b1; // Expected: {'sum': 77, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b10001111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1959,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 77, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001111; b = 8'b11101010; cin = 1'b0; // Expected: {'sum': 57, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001111; b = 8'b11101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1960,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 57, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001100; b = 8'b00000100; cin = 1'b1; // Expected: {'sum': 17, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001100; b = 8'b00000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1961,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 17, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b10001010; cin = 1'b1; // Expected: {'sum': 90, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b10001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1962,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 90, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b00000111; cin = 1'b1; // Expected: {'sum': 147, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b00000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1963,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 147, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b10010110; cin = 1'b1; // Expected: {'sum': 180, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b10010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1964,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 180, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b10001001; cin = 1'b1; // Expected: {'sum': 45, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b10001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1965,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 45, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b01110010; cin = 1'b0; // Expected: {'sum': 142, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b01110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1966,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 142, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b01010101; cin = 1'b1; // Expected: {'sum': 47, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b01010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1967,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 47, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b11101101; cin = 1'b0; // Expected: {'sum': 115, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b11101101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1968,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 115, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b00111100; cin = 1'b1; // Expected: {'sum': 84, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b00111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1969,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 84, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b01000001; cin = 1'b1; // Expected: {'sum': 205, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b01000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1970,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 205, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b00001100; cin = 1'b0; // Expected: {'sum': 254, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b00001100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1971,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 254, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b01011111; cin = 1'b0; // Expected: {'sum': 105, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b01011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1972,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 105, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101101; b = 8'b10000000; cin = 1'b0; // Expected: {'sum': 45, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101101; b = 8'b10000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1973,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 45, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010101; b = 8'b11001100; cin = 1'b0; // Expected: {'sum': 33, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010101; b = 8'b11001100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1974,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 33, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b01010000; cin = 1'b1; // Expected: {'sum': 80, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b01010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1975,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 80, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010011; b = 8'b10111100; cin = 1'b1; // Expected: {'sum': 16, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010011; b = 8'b10111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1976,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 16, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b01111011; cin = 1'b0; // Expected: {'sum': 167, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b01111011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1977,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 167, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100110; b = 8'b10110011; cin = 1'b1; // Expected: {'sum': 154, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100110; b = 8'b10110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1978,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 154, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111110; b = 8'b01000111; cin = 1'b1; // Expected: {'sum': 134, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111110; b = 8'b01000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1979,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 134, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001001; b = 8'b11101011; cin = 1'b1; // Expected: {'sum': 53, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001001; b = 8'b11101011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1980,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 53, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b00100000; cin = 1'b0; // Expected: {'sum': 56, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b00100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1981,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 56, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b11010001; cin = 1'b0; // Expected: {'sum': 24, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b11010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1982,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 24, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011000; b = 8'b11011000; cin = 1'b0; // Expected: {'sum': 48, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011000; b = 8'b11011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1983,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 48, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b00110010; cin = 1'b0; // Expected: {'sum': 101, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b00110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1984,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 101, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111110; b = 8'b01100000; cin = 1'b1; // Expected: {'sum': 159, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111110; b = 8'b01100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1985,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 159, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011001; b = 8'b01000111; cin = 1'b0; // Expected: {'sum': 96, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011001; b = 8'b01000111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1986,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 96, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000110; b = 8'b11000110; cin = 1'b0; // Expected: {'sum': 140, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000110; b = 8'b11000110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1987,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 140, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111010; b = 8'b00111111; cin = 1'b1; // Expected: {'sum': 58, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111010; b = 8'b00111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1988,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 58, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b10101001; cin = 1'b1; // Expected: {'sum': 234, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b10101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1989,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 234, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001100; b = 8'b01001000; cin = 1'b0; // Expected: {'sum': 212, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001100; b = 8'b01001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1990,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 212, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011000; b = 8'b10110010; cin = 1'b0; // Expected: {'sum': 10, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011000; b = 8'b10110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1991,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000111; b = 8'b00001000; cin = 1'b1; // Expected: {'sum': 208, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000111; b = 8'b00001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1992,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 208, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001001; b = 8'b00100111; cin = 1'b1; // Expected: {'sum': 241, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001001; b = 8'b00100111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1993,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 241, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b01100110; cin = 1'b0; // Expected: {'sum': 229, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b01100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1994,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 229, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011010; b = 8'b01011111; cin = 1'b0; // Expected: {'sum': 57, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011010; b = 8'b01011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1995,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 57, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b11011101; cin = 1'b1; // Expected: {'sum': 126, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b11011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1996,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 126, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b10000110; cin = 1'b1; // Expected: {'sum': 245, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b10000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1997,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 245, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b10110100; cin = 1'b1; // Expected: {'sum': 186, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b10110100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1998,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 186, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b11001010; cin = 1'b0; // Expected: {'sum': 156, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b11001010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1999,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 156, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b01010000; cin = 1'b1; // Expected: {'sum': 50, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b01010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2000,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 50, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b10010101; cin = 1'b1; // Expected: {'sum': 136, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b10010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2001,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 136, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b01100011; cin = 1'b0; // Expected: {'sum': 130, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b01100011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2002,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 130, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b10011100; cin = 1'b1; // Expected: {'sum': 114, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b10011100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2003,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 114, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b11101101; cin = 1'b1; // Expected: {'sum': 184, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b11101101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2004,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 184, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b01100010; cin = 1'b0; // Expected: {'sum': 117, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b01100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2005,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 117, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111000; b = 8'b01111000; cin = 1'b0; // Expected: {'sum': 176, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111000; b = 8'b01111000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2006,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 176, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b10000110; cin = 1'b1; // Expected: {'sum': 116, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b10000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2007,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 116, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110001; b = 8'b10000011; cin = 1'b1; // Expected: {'sum': 181, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110001; b = 8'b10000011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2008,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 181, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001101; b = 8'b11001011; cin = 1'b1; // Expected: {'sum': 217, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001101; b = 8'b11001011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2009,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 217, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100010; b = 8'b01001011; cin = 1'b1; // Expected: {'sum': 46, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100010; b = 8'b01001011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2010,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 46, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b01011111; cin = 1'b1; // Expected: {'sum': 11, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b01011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2011,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 11, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b01101100; cin = 1'b0; // Expected: {'sum': 229, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b01101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2012,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 229, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b11000111; cin = 1'b0; // Expected: {'sum': 209, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b11000111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2013,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 209, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110001; b = 8'b00100001; cin = 1'b0; // Expected: {'sum': 82, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110001; b = 8'b00100001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2014,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 82, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b11011011; cin = 1'b0; // Expected: {'sum': 94, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b11011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2015,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 94, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b01101010; cin = 1'b1; // Expected: {'sum': 0, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b01101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2016,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b10111101; cin = 1'b1; // Expected: {'sum': 99, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b10111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2017,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 99, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b10101001; cin = 1'b1; // Expected: {'sum': 179, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b10101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2018,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 179, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b01001000; cin = 1'b1; // Expected: {'sum': 249, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b01001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2019,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 249, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b11010001; cin = 1'b1; // Expected: {'sum': 136, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b11010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2020,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 136, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011101; b = 8'b01000100; cin = 1'b1; // Expected: {'sum': 34, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011101; b = 8'b01000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2021,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 34, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010101; b = 8'b00011011; cin = 1'b0; // Expected: {'sum': 112, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010101; b = 8'b00011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2022,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 112, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b01010001; cin = 1'b0; // Expected: {'sum': 116, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b01010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2023,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 116, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b00100110; cin = 1'b1; // Expected: {'sum': 62, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b00100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2024,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 62, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b00010000; cin = 1'b0; // Expected: {'sum': 53, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b00010000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2025,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 53, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b11111111; cin = 1'b0; // Expected: {'sum': 157, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b11111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2026,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 157, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b10100000; cin = 1'b1; // Expected: {'sum': 211, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b10100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2027,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 211, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b11100010; cin = 1'b0; // Expected: {'sum': 214, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b11100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2028,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 214, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b10110110; cin = 1'b0; // Expected: {'sum': 145, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b10110110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2029,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 145, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b00111100; cin = 1'b1; // Expected: {'sum': 56, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b00111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2030,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 56, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b10110100; cin = 1'b1; // Expected: {'sum': 71, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b10110100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2031,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 71, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b10011100; cin = 1'b1; // Expected: {'sum': 59, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b10011100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2032,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 59, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011001; b = 8'b11011110; cin = 1'b1; // Expected: {'sum': 56, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011001; b = 8'b11011110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2033,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 56, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000001; b = 8'b01001101; cin = 1'b0; // Expected: {'sum': 14, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000001; b = 8'b01001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2034,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101010; b = 8'b11111010; cin = 1'b1; // Expected: {'sum': 229, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101010; b = 8'b11111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2035,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 229, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b01011110; cin = 1'b1; // Expected: {'sum': 145, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b01011110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2036,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 145, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100111; b = 8'b01110000; cin = 1'b0; // Expected: {'sum': 215, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100111; b = 8'b01110000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2037,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 215, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b00111110; cin = 1'b1; // Expected: {'sum': 246, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b00111110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2038,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 246, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b01010110; cin = 1'b0; // Expected: {'sum': 183, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b01010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2039,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 183, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b01110001; cin = 1'b0; // Expected: {'sum': 121, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b01110001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2040,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 121, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b01010011; cin = 1'b0; // Expected: {'sum': 160, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b01010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2041,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 160, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011001; b = 8'b00010100; cin = 1'b1; // Expected: {'sum': 110, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011001; b = 8'b00010100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2042,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 110, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b11011011; cin = 1'b1; // Expected: {'sum': 251, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b11011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2043,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 251, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b01000011; cin = 1'b1; // Expected: {'sum': 91, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b01000011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2044,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 91, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b10000010; cin = 1'b1; // Expected: {'sum': 43, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b10000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2045,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 43, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101010; b = 8'b11011010; cin = 1'b0; // Expected: {'sum': 196, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101010; b = 8'b11011010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2046,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 196, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011110; b = 8'b11111000; cin = 1'b0; // Expected: {'sum': 214, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011110; b = 8'b11111000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2047,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 214, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101011; b = 8'b11001111; cin = 1'b0; // Expected: {'sum': 250, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101011; b = 8'b11001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2048,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 250, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b01000001; cin = 1'b0; // Expected: {'sum': 199, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b01000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2049,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 199, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b10000110; cin = 1'b1; // Expected: {'sum': 144, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b10000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2050,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 144, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b01100101; cin = 1'b1; // Expected: {'sum': 11, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b01100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2051,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 11, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010110; b = 8'b10000110; cin = 1'b1; // Expected: {'sum': 93, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010110; b = 8'b10000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2052,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 93, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b10110000; cin = 1'b1; // Expected: {'sum': 140, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b10110000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2053,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 140, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110001; b = 8'b00100110; cin = 1'b1; // Expected: {'sum': 152, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110001; b = 8'b00100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2054,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 152, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b00001001; cin = 1'b1; // Expected: {'sum': 190, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b00001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2055,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 190, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000011; b = 8'b10110011; cin = 1'b1; // Expected: {'sum': 119, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000011; b = 8'b10110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2056,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 119, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b10001010; cin = 1'b0; // Expected: {'sum': 97, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b10001010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2057,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 97, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b01000111; cin = 1'b0; // Expected: {'sum': 21, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b01000111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2058,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 21, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b10110010; cin = 1'b1; // Expected: {'sum': 47, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b10110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2059,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 47, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b01100011; cin = 1'b0; // Expected: {'sum': 159, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b01100011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2060,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 159, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b00010101; cin = 1'b1; // Expected: {'sum': 3, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b00010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2061,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110111; b = 8'b10110110; cin = 1'b0; // Expected: {'sum': 237, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110111; b = 8'b10110110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2062,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 237, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b00001000; cin = 1'b0; // Expected: {'sum': 76, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b00001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2063,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 76, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010100; b = 8'b11111101; cin = 1'b1; // Expected: {'sum': 18, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010100; b = 8'b11111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2064,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 18, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b00010111; cin = 1'b0; // Expected: {'sum': 14, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b00010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2065,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b10110011; cin = 1'b0; // Expected: {'sum': 42, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b10110011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2066,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 42, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b11111011; cin = 1'b1; // Expected: {'sum': 31, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b11111011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2067,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 31, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101001; b = 8'b10101000; cin = 1'b0; // Expected: {'sum': 17, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101001; b = 8'b10101000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2068,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 17, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011110; b = 8'b00101100; cin = 1'b0; // Expected: {'sum': 10, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011110; b = 8'b00101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2069,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000001; b = 8'b10010010; cin = 1'b0; // Expected: {'sum': 83, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000001; b = 8'b10010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2070,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 83, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001000; b = 8'b11110000; cin = 1'b0; // Expected: {'sum': 56, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001000; b = 8'b11110000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2071,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 56, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b11111001; cin = 1'b1; // Expected: {'sum': 179, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b11111001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2072,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 179, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b00010011; cin = 1'b1; // Expected: {'sum': 111, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b00010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2073,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 111, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b10011111; cin = 1'b0; // Expected: {'sum': 168, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b10011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2074,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 168, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b01110100; cin = 1'b1; // Expected: {'sum': 143, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b01110100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2075,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 143, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100000; b = 8'b11101000; cin = 1'b0; // Expected: {'sum': 72, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100000; b = 8'b11101000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2076,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 72, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b01001011; cin = 1'b0; // Expected: {'sum': 3, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b01001011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2077,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b10111010; cin = 1'b0; // Expected: {'sum': 85, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b10111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2078,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 85, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b10001110; cin = 1'b1; // Expected: {'sum': 7, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b10001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2079,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110100; b = 8'b10100110; cin = 1'b1; // Expected: {'sum': 27, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110100; b = 8'b10100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2080,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 27, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b11000110; cin = 1'b1; // Expected: {'sum': 229, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b11000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2081,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 229, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b00010100; cin = 1'b1; // Expected: {'sum': 213, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b00010100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2082,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 213, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b10110110; cin = 1'b1; // Expected: {'sum': 110, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b10110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2083,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 110, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b00111011; cin = 1'b0; // Expected: {'sum': 198, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b00111011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2084,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 198, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b11011100; cin = 1'b1; // Expected: {'sum': 231, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b11011100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2085,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 231, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010011; b = 8'b11110000; cin = 1'b1; // Expected: {'sum': 196, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010011; b = 8'b11110000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2086,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 196, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b01000111; cin = 1'b1; // Expected: {'sum': 136, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b01000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2087,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 136, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100111; b = 8'b10101101; cin = 1'b1; // Expected: {'sum': 21, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100111; b = 8'b10101101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2088,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 21, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b10111101; cin = 1'b0; // Expected: {'sum': 170, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b10111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2089,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 170, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b00011101; cin = 1'b0; // Expected: {'sum': 38, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b00011101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2090,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 38, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011001; b = 8'b11000111; cin = 1'b1; // Expected: {'sum': 97, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011001; b = 8'b11000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2091,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 97, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111001; b = 8'b11001101; cin = 1'b1; // Expected: {'sum': 7, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111001; b = 8'b11001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2092,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b11010010; cin = 1'b0; // Expected: {'sum': 53, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b11010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2093,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 53, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b01111101; cin = 1'b0; // Expected: {'sum': 189, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b01111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2094,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 189, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111010; b = 8'b10110011; cin = 1'b0; // Expected: {'sum': 173, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111010; b = 8'b10110011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2095,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 173, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b01010111; cin = 1'b1; // Expected: {'sum': 49, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b01010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2096,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 49, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110000; b = 8'b10101111; cin = 1'b1; // Expected: {'sum': 32, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110000; b = 8'b10101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2097,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 32, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100000; b = 8'b10010010; cin = 1'b1; // Expected: {'sum': 115, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100000; b = 8'b10010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2098,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 115, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b00001000; cin = 1'b0; // Expected: {'sum': 240, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b00001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2099,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 240, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b00110001; cin = 1'b1; // Expected: {'sum': 195, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b00110001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2100,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 195, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001011; b = 8'b00001000; cin = 1'b0; // Expected: {'sum': 211, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001011; b = 8'b00001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2101,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 211, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b01001001; cin = 1'b0; // Expected: {'sum': 19, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b01001001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2102,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 19, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b11001100; cin = 1'b1; // Expected: {'sum': 200, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b11001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2103,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 200, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010001; b = 8'b01110101; cin = 1'b1; // Expected: {'sum': 71, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010001; b = 8'b01110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2104,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 71, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010100; b = 8'b01011001; cin = 1'b1; // Expected: {'sum': 110, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010100; b = 8'b01011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2105,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 110, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b01100110; cin = 1'b1; // Expected: {'sum': 202, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b01100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2106,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 202, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b10110001; cin = 1'b0; // Expected: {'sum': 82, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b10110001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2107,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 82, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b11101010; cin = 1'b0; // Expected: {'sum': 172, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b11101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2108,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 172, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b11010010; cin = 1'b0; // Expected: {'sum': 14, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b11010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2109,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b00100000; cin = 1'b1; // Expected: {'sum': 222, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b00100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2110,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 222, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b01000000; cin = 1'b1; // Expected: {'sum': 194, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b01000000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2111,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 194, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100111; b = 8'b11001110; cin = 1'b0; // Expected: {'sum': 117, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100111; b = 8'b11001110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2112,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 117, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100110; b = 8'b10101110; cin = 1'b0; // Expected: {'sum': 148, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100110; b = 8'b10101110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2113,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 148, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b11100010; cin = 1'b0; // Expected: {'sum': 193, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b11100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2114,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 193, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b10111001; cin = 1'b0; // Expected: {'sum': 39, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b10111001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2115,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 39, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b10101011; cin = 1'b0; // Expected: {'sum': 121, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b10101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2116,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 121, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b01011111; cin = 1'b0; // Expected: {'sum': 175, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b01011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2117,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 175, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001111; b = 8'b11011011; cin = 1'b0; // Expected: {'sum': 42, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001111; b = 8'b11011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2118,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 42, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b10010110; cin = 1'b1; // Expected: {'sum': 248, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b10010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2119,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 248, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111000; b = 8'b01110110; cin = 1'b1; // Expected: {'sum': 111, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111000; b = 8'b01110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2120,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 111, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b01111011; cin = 1'b1; // Expected: {'sum': 109, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b01111011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2121,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 109, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b11100001; cin = 1'b1; // Expected: {'sum': 219, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b11100001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2122,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 219, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001111; b = 8'b11110101; cin = 1'b0; // Expected: {'sum': 68, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001111; b = 8'b11110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2123,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 68, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b00001000; cin = 1'b0; // Expected: {'sum': 233, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b00001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2124,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 233, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b00011101; cin = 1'b1; // Expected: {'sum': 21, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b00011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2125,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 21, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b00100100; cin = 1'b1; // Expected: {'sum': 46, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b00100100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2126,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 46, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110001; b = 8'b10111100; cin = 1'b0; // Expected: {'sum': 45, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110001; b = 8'b10111100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2127,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 45, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b10001000; cin = 1'b0; // Expected: {'sum': 99, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b10001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2128,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 99, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b00011111; cin = 1'b0; // Expected: {'sum': 135, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b00011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2129,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 135, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b11011011; cin = 1'b1; // Expected: {'sum': 32, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b11011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2130,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 32, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b10010010; cin = 1'b1; // Expected: {'sum': 181, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b10010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2131,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 181, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b10011000; cin = 1'b0; // Expected: {'sum': 81, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b10011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2132,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 81, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b10100011; cin = 1'b0; // Expected: {'sum': 14, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b10100011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2133,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b11100111; cin = 1'b1; // Expected: {'sum': 219, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b11100111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2134,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 219, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b10101101; cin = 1'b0; // Expected: {'sum': 66, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b10101101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2135,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 66, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b00000110; cin = 1'b0; // Expected: {'sum': 15, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b00000110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2136,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b00101000; cin = 1'b0; // Expected: {'sum': 148, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b00101000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2137,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 148, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b01010011; cin = 1'b0; // Expected: {'sum': 193, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b01010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2138,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 193, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111011; b = 8'b11001111; cin = 1'b0; // Expected: {'sum': 10, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111011; b = 8'b11001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2139,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001001; b = 8'b11100010; cin = 1'b0; // Expected: {'sum': 171, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001001; b = 8'b11100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2140,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 171, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b01101011; cin = 1'b0; // Expected: {'sum': 70, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b01101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2141,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 70, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010011; b = 8'b00001011; cin = 1'b0; // Expected: {'sum': 222, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010011; b = 8'b00001011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2142,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 222, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b10101001; cin = 1'b0; // Expected: {'sum': 12, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b10101001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2143,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b11100100; cin = 1'b1; // Expected: {'sum': 165, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b11100100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2144,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 165, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b00110010; cin = 1'b0; // Expected: {'sum': 165, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b00110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2145,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 165, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010111; b = 8'b10110010; cin = 1'b0; // Expected: {'sum': 9, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010111; b = 8'b10110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2146,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 9, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010110; b = 8'b01100101; cin = 1'b0; // Expected: {'sum': 59, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010110; b = 8'b01100101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2147,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 59, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b11111111; cin = 1'b1; // Expected: {'sum': 246, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b11111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2148,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 246, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b00101100; cin = 1'b0; // Expected: {'sum': 3, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b00101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2149,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011011; b = 8'b01111000; cin = 1'b0; // Expected: {'sum': 147, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011011; b = 8'b01111000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2150,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 147, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011101; b = 8'b11010010; cin = 1'b0; // Expected: {'sum': 111, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011101; b = 8'b11010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2151,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 111, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b00010011; cin = 1'b0; // Expected: {'sum': 169, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b00010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2152,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 169, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b01110101; cin = 1'b1; // Expected: {'sum': 111, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b01110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2153,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 111, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b00011100; cin = 1'b1; // Expected: {'sum': 126, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b00011100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2154,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 126, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111011; b = 8'b11111010; cin = 1'b0; // Expected: {'sum': 181, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111011; b = 8'b11111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2155,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 181, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101010; b = 8'b00010111; cin = 1'b1; // Expected: {'sum': 194, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101010; b = 8'b00010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2156,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 194, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b01101101; cin = 1'b0; // Expected: {'sum': 233, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b01101101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2157,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 233, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000110; b = 8'b00100010; cin = 1'b0; // Expected: {'sum': 40, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000110; b = 8'b00100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2158,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 40, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b11011011; cin = 1'b0; // Expected: {'sum': 40, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b11011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2159,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 40, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b10000010; cin = 1'b0; // Expected: {'sum': 245, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b10000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2160,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 245, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b01111101; cin = 1'b0; // Expected: {'sum': 86, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b01111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2161,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 86, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b01111001; cin = 1'b0; // Expected: {'sum': 221, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b01111001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2162,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 221, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b11100011; cin = 1'b0; // Expected: {'sum': 90, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b11100011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2163,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 90, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b01111101; cin = 1'b0; // Expected: {'sum': 206, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b01111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2164,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 206, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b11011101; cin = 1'b1; // Expected: {'sum': 156, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b11011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2165,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 156, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b00000001; cin = 1'b0; // Expected: {'sum': 151, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b00000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2166,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 151, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b01001100; cin = 1'b0; // Expected: {'sum': 167, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b01001100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2167,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 167, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b10110100; cin = 1'b0; // Expected: {'sum': 120, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b10110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2168,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 120, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010111; b = 8'b10011010; cin = 1'b1; // Expected: {'sum': 242, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010111; b = 8'b10011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2169,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 242, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100010; b = 8'b10001010; cin = 1'b1; // Expected: {'sum': 45, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100010; b = 8'b10001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2170,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 45, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b10011000; cin = 1'b0; // Expected: {'sum': 145, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b10011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2171,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 145, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b00100101; cin = 1'b1; // Expected: {'sum': 213, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b00100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2172,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 213, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110001; b = 8'b11000001; cin = 1'b1; // Expected: {'sum': 51, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110001; b = 8'b11000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2173,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 51, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b01110010; cin = 1'b1; // Expected: {'sum': 213, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b01110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2174,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 213, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011111; b = 8'b01101001; cin = 1'b1; // Expected: {'sum': 201, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011111; b = 8'b01101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2175,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 201, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b01101110; cin = 1'b0; // Expected: {'sum': 217, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b01101110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2176,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 217, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001000; b = 8'b11100110; cin = 1'b0; // Expected: {'sum': 174, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001000; b = 8'b11100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2177,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 174, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b10101110; cin = 1'b1; // Expected: {'sum': 5, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b10101110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2178,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 5, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b01001111; cin = 1'b0; // Expected: {'sum': 11, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b01001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2179,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 11, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b00011111; cin = 1'b0; // Expected: {'sum': 146, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b00011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2180,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 146, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b11010001; cin = 1'b1; // Expected: {'sum': 109, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b11010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2181,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 109, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b01110101; cin = 1'b1; // Expected: {'sum': 149, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b01110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2182,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 149, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b11011010; cin = 1'b1; // Expected: {'sum': 215, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b11011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2183,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 215, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b11100101; cin = 1'b1; // Expected: {'sum': 0, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b11100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2184,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111011; b = 8'b00000010; cin = 1'b1; // Expected: {'sum': 126, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111011; b = 8'b00000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2185,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 126, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b10010111; cin = 1'b1; // Expected: {'sum': 51, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b10010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2186,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 51, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b10001000; cin = 1'b0; // Expected: {'sum': 62, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b10001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2187,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 62, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b01000100; cin = 1'b0; // Expected: {'sum': 54, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b01000100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2188,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 54, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b00000110; cin = 1'b1; // Expected: {'sum': 132, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b00000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2189,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 132, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b01010001; cin = 1'b0; // Expected: {'sum': 81, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b01010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2190,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 81, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b10001111; cin = 1'b1; // Expected: {'sum': 40, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b10001111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2191,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 40, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b10010010; cin = 1'b1; // Expected: {'sum': 74, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b10010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2192,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 74, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011000; b = 8'b11000011; cin = 1'b0; // Expected: {'sum': 27, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011000; b = 8'b11000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2193,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 27, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b10101001; cin = 1'b1; // Expected: {'sum': 152, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b10101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2194,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 152, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b11001110; cin = 1'b0; // Expected: {'sum': 92, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b11001110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2195,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 92, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b11001000; cin = 1'b0; // Expected: {'sum': 190, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b11001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2196,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 190, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011111; b = 8'b01100110; cin = 1'b1; // Expected: {'sum': 198, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011111; b = 8'b01100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2197,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 198, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b10011011; cin = 1'b1; // Expected: {'sum': 63, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b10011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2198,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 63, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111111; b = 8'b00001101; cin = 1'b0; // Expected: {'sum': 204, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111111; b = 8'b00001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2199,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 204, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b10100011; cin = 1'b1; // Expected: {'sum': 188, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b10100011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2200,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 188, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b11011101; cin = 1'b0; // Expected: {'sum': 99, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b11011101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2201,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 99, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001011; b = 8'b00000111; cin = 1'b0; // Expected: {'sum': 18, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001011; b = 8'b00000111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2202,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 18, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b11011001; cin = 1'b0; // Expected: {'sum': 206, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b11011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2203,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 206, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b01101111; cin = 1'b1; // Expected: {'sum': 140, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b01101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2204,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 140, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b01111000; cin = 1'b0; // Expected: {'sum': 128, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b01111000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2205,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 128, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111101; b = 8'b11110000; cin = 1'b1; // Expected: {'sum': 238, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111101; b = 8'b11110000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2206,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 238, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b11010001; cin = 1'b0; // Expected: {'sum': 103, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b11010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2207,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 103, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b10000110; cin = 1'b1; // Expected: {'sum': 123, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b10000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2208,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 123, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b01001101; cin = 1'b0; // Expected: {'sum': 118, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b01001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2209,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 118, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b00110101; cin = 1'b0; // Expected: {'sum': 134, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b00110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2210,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 134, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b00101111; cin = 1'b1; // Expected: {'sum': 145, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b00101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2211,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 145, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b10010111; cin = 1'b0; // Expected: {'sum': 144, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b10010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2212,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 144, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b11101110; cin = 1'b1; // Expected: {'sum': 158, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b11101110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2213,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 158, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b10010000; cin = 1'b1; // Expected: {'sum': 114, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b10010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2214,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 114, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010100; b = 8'b01011101; cin = 1'b1; // Expected: {'sum': 114, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010100; b = 8'b01011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2215,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 114, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b00000101; cin = 1'b1; // Expected: {'sum': 135, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b00000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2216,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 135, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001101; b = 8'b11011100; cin = 1'b1; // Expected: {'sum': 234, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001101; b = 8'b11011100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2217,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 234, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b01100101; cin = 1'b0; // Expected: {'sum': 99, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b01100101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2218,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 99, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010011; b = 8'b10011011; cin = 1'b0; // Expected: {'sum': 110, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010011; b = 8'b10011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2219,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 110, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b11110000; cin = 1'b0; // Expected: {'sum': 114, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b11110000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2220,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 114, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010100; b = 8'b00001110; cin = 1'b0; // Expected: {'sum': 34, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010100; b = 8'b00001110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2221,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 34, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010001; b = 8'b11111111; cin = 1'b0; // Expected: {'sum': 208, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010001; b = 8'b11111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2222,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 208, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b01011010; cin = 1'b1; // Expected: {'sum': 149, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b01011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2223,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 149, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b11111111; cin = 1'b0; // Expected: {'sum': 140, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b11111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2224,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 140, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b01011011; cin = 1'b1; // Expected: {'sum': 142, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b01011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2225,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 142, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110110; b = 8'b01110101; cin = 1'b0; // Expected: {'sum': 235, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110110; b = 8'b01110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2226,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 235, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b10111000; cin = 1'b1; // Expected: {'sum': 75, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b10111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2227,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 75, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100100; b = 8'b00101111; cin = 1'b0; // Expected: {'sum': 211, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100100; b = 8'b00101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2228,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 211, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111111; b = 8'b11100000; cin = 1'b1; // Expected: {'sum': 32, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111111; b = 8'b11100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2229,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 32, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b10110100; cin = 1'b1; // Expected: {'sum': 188, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b10110100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2230,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 188, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100110; b = 8'b00001101; cin = 1'b0; // Expected: {'sum': 243, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100110; b = 8'b00001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2231,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 243, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101001; b = 8'b00001010; cin = 1'b1; // Expected: {'sum': 244, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101001; b = 8'b00001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2232,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 244, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b01011011; cin = 1'b0; // Expected: {'sum': 101, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b01011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2233,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 101, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b00111100; cin = 1'b1; // Expected: {'sum': 96, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b00111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2234,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 96, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b10101100; cin = 1'b1; // Expected: {'sum': 125, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b10101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2235,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 125, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110001; b = 8'b11000110; cin = 1'b1; // Expected: {'sum': 248, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110001; b = 8'b11000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2236,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 248, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b10110011; cin = 1'b1; // Expected: {'sum': 188, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b10110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2237,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 188, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b11001110; cin = 1'b1; // Expected: {'sum': 191, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b11001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2238,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 191, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b00000010; cin = 1'b0; // Expected: {'sum': 7, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b00000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2239,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101011; b = 8'b01110100; cin = 1'b0; // Expected: {'sum': 159, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101011; b = 8'b01110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2240,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 159, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b01100001; cin = 1'b0; // Expected: {'sum': 223, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b01100001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2241,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 223, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100110; b = 8'b11011110; cin = 1'b1; // Expected: {'sum': 5, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100110; b = 8'b11011110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2242,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 5, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111111; b = 8'b00101101; cin = 1'b1; // Expected: {'sum': 237, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111111; b = 8'b00101101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2243,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 237, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b00110100; cin = 1'b1; // Expected: {'sum': 190, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b00110100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2244,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 190, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b00111101; cin = 1'b0; // Expected: {'sum': 192, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b00111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2245,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 192, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b00110000; cin = 1'b1; // Expected: {'sum': 204, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b00110000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2246,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 204, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000111; b = 8'b10110001; cin = 1'b1; // Expected: {'sum': 121, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000111; b = 8'b10110001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2247,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 121, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111011; b = 8'b01100100; cin = 1'b1; // Expected: {'sum': 224, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111011; b = 8'b01100100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2248,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 224, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011001; b = 8'b10011101; cin = 1'b1; // Expected: {'sum': 247, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011001; b = 8'b10011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2249,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 247, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111011; b = 8'b01101111; cin = 1'b0; // Expected: {'sum': 170, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111011; b = 8'b01101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2250,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 170, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b00111100; cin = 1'b0; // Expected: {'sum': 153, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b00111100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2251,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 153, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b00010111; cin = 1'b0; // Expected: {'sum': 209, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b00010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2252,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 209, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b10001111; cin = 1'b0; // Expected: {'sum': 8, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b10001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2253,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 8, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b11010001; cin = 1'b0; // Expected: {'sum': 29, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b11010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2254,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 29, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b10010000; cin = 1'b1; // Expected: {'sum': 118, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b10010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2255,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 118, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b01101000; cin = 1'b1; // Expected: {'sum': 39, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b01101000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2256,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 39, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b10111101; cin = 1'b1; // Expected: {'sum': 150, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b10111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2257,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 150, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110010; b = 8'b10101001; cin = 1'b0; // Expected: {'sum': 27, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110010; b = 8'b10101001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2258,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 27, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111110; b = 8'b01000000; cin = 1'b1; // Expected: {'sum': 127, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111110; b = 8'b01000000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2259,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 127, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b00010111; cin = 1'b1; // Expected: {'sum': 167, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b00010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2260,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 167, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b10000011; cin = 1'b0; // Expected: {'sum': 90, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b10000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2261,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 90, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b11011000; cin = 1'b0; // Expected: {'sum': 59, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b11011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2262,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 59, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b11010001; cin = 1'b1; // Expected: {'sum': 98, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b11010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2263,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 98, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b10100000; cin = 1'b0; // Expected: {'sum': 75, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b10100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2264,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 75, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011010; b = 8'b01101001; cin = 1'b1; // Expected: {'sum': 196, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011010; b = 8'b01101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2265,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 196, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010101; b = 8'b01101001; cin = 1'b0; // Expected: {'sum': 126, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010101; b = 8'b01101001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2266,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 126, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b10110110; cin = 1'b0; // Expected: {'sum': 134, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b10110110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2267,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 134, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b01110011; cin = 1'b0; // Expected: {'sum': 191, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b01110011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2268,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 191, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b11111011; cin = 1'b0; // Expected: {'sum': 93, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b11111011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2269,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 93, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b11000011; cin = 1'b0; // Expected: {'sum': 194, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b11000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2270,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 194, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b10010111; cin = 1'b0; // Expected: {'sum': 187, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b10010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2271,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 187, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b10000101; cin = 1'b0; // Expected: {'sum': 90, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b10000101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2272,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 90, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b10011111; cin = 1'b0; // Expected: {'sum': 119, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b10011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2273,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 119, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b11000111; cin = 1'b1; // Expected: {'sum': 152, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b11000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2274,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 152, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b00101001; cin = 1'b0; // Expected: {'sum': 196, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b00101001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2275,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 196, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100100; b = 8'b00010110; cin = 1'b0; // Expected: {'sum': 186, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100100; b = 8'b00010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2276,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 186, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b11010010; cin = 1'b0; // Expected: {'sum': 64, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b11010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2277,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 64, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b01101001; cin = 1'b1; // Expected: {'sum': 238, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b01101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2278,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 238, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111111; b = 8'b11110101; cin = 1'b1; // Expected: {'sum': 181, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111111; b = 8'b11110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2279,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 181, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b00001101; cin = 1'b0; // Expected: {'sum': 226, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b00001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2280,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 226, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101111; b = 8'b10101001; cin = 1'b1; // Expected: {'sum': 217, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101111; b = 8'b10101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2281,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 217, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b00110010; cin = 1'b1; // Expected: {'sum': 115, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b00110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2282,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 115, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100111; b = 8'b10110100; cin = 1'b1; // Expected: {'sum': 156, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100111; b = 8'b10110100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2283,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 156, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b01101000; cin = 1'b0; // Expected: {'sum': 61, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b01101000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2284,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 61, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b01101101; cin = 1'b0; // Expected: {'sum': 224, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b01101101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2285,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 224, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b11000000; cin = 1'b1; // Expected: {'sum': 238, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b11000000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2286,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 238, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b11011110; cin = 1'b0; // Expected: {'sum': 208, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b11011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2287,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 208, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110100; b = 8'b10111010; cin = 1'b0; // Expected: {'sum': 46, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110100; b = 8'b10111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2288,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 46, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b10100111; cin = 1'b0; // Expected: {'sum': 243, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b10100111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2289,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 243, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111011; b = 8'b01101111; cin = 1'b1; // Expected: {'sum': 43, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111011; b = 8'b01101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2290,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 43, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100110; b = 8'b11001011; cin = 1'b0; // Expected: {'sum': 241, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100110; b = 8'b11001011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2291,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 241, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b10100110; cin = 1'b0; // Expected: {'sum': 42, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b10100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2292,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 42, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100010; b = 8'b00100010; cin = 1'b1; // Expected: {'sum': 197, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100010; b = 8'b00100010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2293,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 197, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b10000000; cin = 1'b0; // Expected: {'sum': 58, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b10000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2294,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 58, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010110; b = 8'b11111001; cin = 1'b1; // Expected: {'sum': 208, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010110; b = 8'b11111001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2295,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 208, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b01001000; cin = 1'b0; // Expected: {'sum': 222, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b01001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2296,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 222, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100100; b = 8'b01010000; cin = 1'b0; // Expected: {'sum': 244, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100100; b = 8'b01010000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2297,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 244, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b11011010; cin = 1'b1; // Expected: {'sum': 92, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b11011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2298,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 92, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100001; b = 8'b01010010; cin = 1'b0; // Expected: {'sum': 115, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100001; b = 8'b01010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2299,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 115, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b11011111; cin = 1'b1; // Expected: {'sum': 229, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b11011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2300,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 229, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b10101111; cin = 1'b1; // Expected: {'sum': 193, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b10101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2301,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 193, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011001; b = 8'b11100101; cin = 1'b1; // Expected: {'sum': 127, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011001; b = 8'b11100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2302,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 127, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b11001110; cin = 1'b0; // Expected: {'sum': 89, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b11001110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2303,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 89, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b00111111; cin = 1'b0; // Expected: {'sum': 71, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b00111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2304,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 71, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b11101010; cin = 1'b1; // Expected: {'sum': 130, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b11101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2305,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 130, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b11110101; cin = 1'b0; // Expected: {'sum': 173, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b11110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2306,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 173, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100111; b = 8'b10001101; cin = 1'b0; // Expected: {'sum': 244, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100111; b = 8'b10001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2307,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 244, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b00101010; cin = 1'b1; // Expected: {'sum': 186, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b00101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2308,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 186, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100110; b = 8'b10101011; cin = 1'b0; // Expected: {'sum': 145, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100110; b = 8'b10101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2309,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 145, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b10101100; cin = 1'b0; // Expected: {'sum': 48, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b10101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2310,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 48, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b11001111; cin = 1'b0; // Expected: {'sum': 197, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b11001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2311,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 197, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b01001111; cin = 1'b1; // Expected: {'sum': 212, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b01001111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2312,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 212, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b11110001; cin = 1'b0; // Expected: {'sum': 242, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b11110001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2313,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 242, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010100; b = 8'b00100101; cin = 1'b1; // Expected: {'sum': 186, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010100; b = 8'b00100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2314,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 186, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b01010110; cin = 1'b0; // Expected: {'sum': 232, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b01010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2315,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 232, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100001; b = 8'b10100111; cin = 1'b1; // Expected: {'sum': 201, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100001; b = 8'b10100111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2316,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 201, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001010; b = 8'b11100011; cin = 1'b1; // Expected: {'sum': 110, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001010; b = 8'b11100011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2317,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 110, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b10001110; cin = 1'b0; // Expected: {'sum': 38, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b10001110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2318,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 38, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b11111101; cin = 1'b1; // Expected: {'sum': 206, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b11111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2319,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 206, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110101; b = 8'b11000010; cin = 1'b0; // Expected: {'sum': 247, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110101; b = 8'b11000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2320,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 247, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b11010111; cin = 1'b1; // Expected: {'sum': 136, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b11010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2321,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 136, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b00010010; cin = 1'b0; // Expected: {'sum': 200, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b00010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2322,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 200, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001000; b = 8'b01110110; cin = 1'b1; // Expected: {'sum': 191, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001000; b = 8'b01110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2323,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 191, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b00000100; cin = 1'b0; // Expected: {'sum': 64, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b00000100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2324,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 64, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b01101101; cin = 1'b0; // Expected: {'sum': 100, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b01101101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2325,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 100, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110111; b = 8'b10111110; cin = 1'b1; // Expected: {'sum': 246, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110111; b = 8'b10111110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2326,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 246, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001111; b = 8'b11111010; cin = 1'b1; // Expected: {'sum': 10, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001111; b = 8'b11111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2327,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b01001111; cin = 1'b1; // Expected: {'sum': 89, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b01001111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2328,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 89, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b00000111; cin = 1'b1; // Expected: {'sum': 53, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b00000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2329,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 53, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b00000011; cin = 1'b0; // Expected: {'sum': 149, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b00000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2330,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 149, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000101; b = 8'b11101000; cin = 1'b1; // Expected: {'sum': 110, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000101; b = 8'b11101000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2331,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 110, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b00010001; cin = 1'b0; // Expected: {'sum': 224, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b00010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2332,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 224, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101100; b = 8'b00111100; cin = 1'b1; // Expected: {'sum': 41, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101100; b = 8'b00111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2333,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 41, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111110; b = 8'b10011011; cin = 1'b0; // Expected: {'sum': 217, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111110; b = 8'b10011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2334,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 217, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110110; b = 8'b00001111; cin = 1'b1; // Expected: {'sum': 134, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110110; b = 8'b00001111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2335,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 134, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b00010010; cin = 1'b1; // Expected: {'sum': 20, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b00010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2336,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 20, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110100; b = 8'b10001000; cin = 1'b0; // Expected: {'sum': 252, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110100; b = 8'b10001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2337,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 252, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b01111010; cin = 1'b1; // Expected: {'sum': 83, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b01111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2338,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 83, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b01101001; cin = 1'b1; // Expected: {'sum': 11, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b01101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2339,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 11, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111111; b = 8'b00001110; cin = 1'b0; // Expected: {'sum': 77, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111111; b = 8'b00001110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2340,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 77, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001101; b = 8'b11010000; cin = 1'b1; // Expected: {'sum': 222, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001101; b = 8'b11010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2341,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 222, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101111; b = 8'b00111110; cin = 1'b0; // Expected: {'sum': 45, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101111; b = 8'b00111110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2342,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 45, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b11010011; cin = 1'b1; // Expected: {'sum': 150, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b11010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2343,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 150, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b10001000; cin = 1'b1; // Expected: {'sum': 83, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b10001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2344,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 83, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b00100110; cin = 1'b1; // Expected: {'sum': 108, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b00100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2345,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 108, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010010; b = 8'b10010001; cin = 1'b0; // Expected: {'sum': 163, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010010; b = 8'b10010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2346,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 163, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110010; b = 8'b01110110; cin = 1'b1; // Expected: {'sum': 233, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110010; b = 8'b01110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2347,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 233, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b11001010; cin = 1'b0; // Expected: {'sum': 20, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b11001010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2348,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 20, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001110; b = 8'b10010010; cin = 1'b1; // Expected: {'sum': 161, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001110; b = 8'b10010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2349,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 161, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b11111111; cin = 1'b0; // Expected: {'sum': 236, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b11111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2350,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 236, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111111; b = 8'b10001001; cin = 1'b1; // Expected: {'sum': 73, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111111; b = 8'b10001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2351,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 73, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111101; b = 8'b00100010; cin = 1'b0; // Expected: {'sum': 31, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111101; b = 8'b00100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2352,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 31, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101001; b = 8'b10000101; cin = 1'b0; // Expected: {'sum': 238, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101001; b = 8'b10000101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2353,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 238, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b01100000; cin = 1'b1; // Expected: {'sum': 163, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b01100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2354,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 163, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b10011111; cin = 1'b1; // Expected: {'sum': 53, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b10011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2355,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 53, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b00001110; cin = 1'b1; // Expected: {'sum': 20, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b00001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2356,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 20, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b11100110; cin = 1'b0; // Expected: {'sum': 93, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b11100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2357,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 93, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b01000110; cin = 1'b0; // Expected: {'sum': 70, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b01000110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2358,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 70, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b11000011; cin = 1'b0; // Expected: {'sum': 38, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b11000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2359,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 38, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b10100000; cin = 1'b1; // Expected: {'sum': 89, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b10100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2360,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 89, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011111; b = 8'b00011110; cin = 1'b0; // Expected: {'sum': 189, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011111; b = 8'b00011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2361,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 189, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100000; b = 8'b01101111; cin = 1'b0; // Expected: {'sum': 79, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100000; b = 8'b01101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2362,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 79, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011001; b = 8'b10001011; cin = 1'b0; // Expected: {'sum': 36, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011001; b = 8'b10001011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2363,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 36, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b10001110; cin = 1'b0; // Expected: {'sum': 193, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b10001110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2364,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 193, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b00000010; cin = 1'b0; // Expected: {'sum': 170, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b00000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2365,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 170, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101100; b = 8'b11110001; cin = 1'b0; // Expected: {'sum': 221, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101100; b = 8'b11110001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2366,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 221, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b00000101; cin = 1'b0; // Expected: {'sum': 222, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b00000101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2367,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 222, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010101; b = 8'b11100110; cin = 1'b0; // Expected: {'sum': 251, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010101; b = 8'b11100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2368,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 251, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b10010110; cin = 1'b1; // Expected: {'sum': 16, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b10010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2369,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 16, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111000; b = 8'b01010001; cin = 1'b0; // Expected: {'sum': 73, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111000; b = 8'b01010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2370,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 73, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b00001111; cin = 1'b0; // Expected: {'sum': 158, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b00001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2371,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 158, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b00001011; cin = 1'b0; // Expected: {'sum': 171, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b00001011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2372,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 171, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b00011011; cin = 1'b0; // Expected: {'sum': 23, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b00011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2373,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 23, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b11110010; cin = 1'b1; // Expected: {'sum': 212, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b11110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2374,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 212, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b00110111; cin = 1'b1; // Expected: {'sum': 183, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b00110111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2375,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 183, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b00011010; cin = 1'b1; // Expected: {'sum': 166, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b00011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2376,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 166, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b01100111; cin = 1'b1; // Expected: {'sum': 40, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b01100111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2377,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 40, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b10010010; cin = 1'b1; // Expected: {'sum': 241, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b10010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2378,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 241, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111111; b = 8'b01000010; cin = 1'b0; // Expected: {'sum': 1, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111111; b = 8'b01000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2379,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b00111111; cin = 1'b1; // Expected: {'sum': 2, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b00111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2380,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b01010110; cin = 1'b0; // Expected: {'sum': 47, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b01010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2381,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 47, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010100; b = 8'b10101000; cin = 1'b1; // Expected: {'sum': 253, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010100; b = 8'b10101000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2382,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 253, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010101; b = 8'b00110100; cin = 1'b1; // Expected: {'sum': 138, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010101; b = 8'b00110100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2383,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 138, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010011; b = 8'b00011110; cin = 1'b0; // Expected: {'sum': 177, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010011; b = 8'b00011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2384,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 177, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b00100000; cin = 1'b1; // Expected: {'sum': 127, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b00100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2385,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 127, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b11010001; cin = 1'b1; // Expected: {'sum': 73, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b11010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2386,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 73, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b10110010; cin = 1'b0; // Expected: {'sum': 16, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b10110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2387,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 16, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011101; b = 8'b01000011; cin = 1'b1; // Expected: {'sum': 33, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011101; b = 8'b01000011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2388,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 33, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b00001000; cin = 1'b0; // Expected: {'sum': 32, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b00001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2389,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 32, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b10111100; cin = 1'b1; // Expected: {'sum': 84, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b10111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2390,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 84, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011001; b = 8'b01111000; cin = 1'b1; // Expected: {'sum': 210, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011001; b = 8'b01111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2391,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 210, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b11011001; cin = 1'b1; // Expected: {'sum': 104, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b11011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2392,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 104, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100010; b = 8'b10000010; cin = 1'b1; // Expected: {'sum': 101, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100010; b = 8'b10000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2393,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 101, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b00111000; cin = 1'b1; // Expected: {'sum': 38, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b00111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2394,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 38, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000011; b = 8'b10100001; cin = 1'b1; // Expected: {'sum': 165, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000011; b = 8'b10100001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2395,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 165, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100111; b = 8'b01110110; cin = 1'b0; // Expected: {'sum': 157, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100111; b = 8'b01110110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2396,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 157, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111000; b = 8'b11000110; cin = 1'b0; // Expected: {'sum': 190, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111000; b = 8'b11000110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2397,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 190, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b11011000; cin = 1'b0; // Expected: {'sum': 214, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b11011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2398,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 214, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b11010110; cin = 1'b1; // Expected: {'sum': 100, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b11010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2399,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 100, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b00100000; cin = 1'b1; // Expected: {'sum': 0, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b00100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2400,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b11111010; cin = 1'b0; // Expected: {'sum': 125, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b11111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2401,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 125, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b00110111; cin = 1'b0; // Expected: {'sum': 106, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b00110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2402,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 106, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b10001001; cin = 1'b0; // Expected: {'sum': 252, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b10001001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2403,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 252, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b10010011; cin = 1'b1; // Expected: {'sum': 33, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b10010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2404,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 33, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111111; b = 8'b11101001; cin = 1'b0; // Expected: {'sum': 168, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111111; b = 8'b11101001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2405,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 168, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001100; b = 8'b00111101; cin = 1'b1; // Expected: {'sum': 74, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001100; b = 8'b00111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2406,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 74, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000100; b = 8'b00010101; cin = 1'b0; // Expected: {'sum': 25, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000100; b = 8'b00010101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2407,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 25, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011001; b = 8'b00000110; cin = 1'b1; // Expected: {'sum': 32, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011001; b = 8'b00000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2408,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 32, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b00010100; cin = 1'b0; // Expected: {'sum': 154, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b00010100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2409,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 154, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b10001111; cin = 1'b0; // Expected: {'sum': 252, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b10001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2410,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 252, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b00000100; cin = 1'b0; // Expected: {'sum': 212, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b00000100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2411,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 212, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b01010011; cin = 1'b1; // Expected: {'sum': 71, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b01010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2412,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 71, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001110; b = 8'b11011001; cin = 1'b1; // Expected: {'sum': 40, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001110; b = 8'b11011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2413,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 40, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101100; b = 8'b10111100; cin = 1'b1; // Expected: {'sum': 105, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101100; b = 8'b10111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2414,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 105, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b00011010; cin = 1'b1; // Expected: {'sum': 177, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b00011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2415,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 177, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011110; b = 8'b11111010; cin = 1'b0; // Expected: {'sum': 216, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011110; b = 8'b11111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2416,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 216, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b11100101; cin = 1'b1; // Expected: {'sum': 68, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b11100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2417,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 68, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b10001110; cin = 1'b1; // Expected: {'sum': 180, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b10001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2418,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 180, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100000; b = 8'b00010000; cin = 1'b1; // Expected: {'sum': 49, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100000; b = 8'b00010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2419,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 49, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b10101110; cin = 1'b0; // Expected: {'sum': 226, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b10101110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2420,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 226, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b10011101; cin = 1'b1; // Expected: {'sum': 157, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b10011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2421,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 157, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b11110100; cin = 1'b0; // Expected: {'sum': 182, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b11110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2422,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 182, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101010; b = 8'b01010111; cin = 1'b0; // Expected: {'sum': 129, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101010; b = 8'b01010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2423,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 129, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011001; b = 8'b00100000; cin = 1'b0; // Expected: {'sum': 57, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011001; b = 8'b00100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2424,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 57, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b11110111; cin = 1'b0; // Expected: {'sum': 100, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b11110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2425,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 100, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b00011100; cin = 1'b1; // Expected: {'sum': 51, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b00011100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2426,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 51, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b00110101; cin = 1'b0; // Expected: {'sum': 120, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b00110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2427,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 120, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b00000000; cin = 1'b0; // Expected: {'sum': 131, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b00000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2428,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 131, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b01001101; cin = 1'b1; // Expected: {'sum': 136, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b01001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2429,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 136, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001111; b = 8'b01110010; cin = 1'b1; // Expected: {'sum': 130, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001111; b = 8'b01110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2430,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 130, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110101; b = 8'b10001011; cin = 1'b0; // Expected: {'sum': 64, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110101; b = 8'b10001011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2431,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 64, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b11000011; cin = 1'b0; // Expected: {'sum': 104, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b11000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2432,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 104, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b01010110; cin = 1'b1; // Expected: {'sum': 156, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b01010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2433,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 156, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b10101001; cin = 1'b1; // Expected: {'sum': 90, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b10101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2434,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 90, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101101; b = 8'b01010110; cin = 1'b0; // Expected: {'sum': 3, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101101; b = 8'b01010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2435,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b10011011; cin = 1'b0; // Expected: {'sum': 148, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b10011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2436,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 148, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b01111001; cin = 1'b1; // Expected: {'sum': 54, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b01111001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2437,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 54, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000100; b = 8'b10001000; cin = 1'b0; // Expected: {'sum': 140, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000100; b = 8'b10001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2438,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 140, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b11100010; cin = 1'b0; // Expected: {'sum': 63, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b11100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2439,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 63, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b11101100; cin = 1'b1; // Expected: {'sum': 100, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b11101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2440,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 100, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001110; b = 8'b10010010; cin = 1'b0; // Expected: {'sum': 224, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001110; b = 8'b10010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2441,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 224, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b11111101; cin = 1'b0; // Expected: {'sum': 74, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b11111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2442,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 74, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b00010001; cin = 1'b0; // Expected: {'sum': 207, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b00010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2443,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 207, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b00001110; cin = 1'b1; // Expected: {'sum': 204, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b00001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2444,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 204, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b11101110; cin = 1'b0; // Expected: {'sum': 131, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b11101110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2445,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 131, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b01001011; cin = 1'b0; // Expected: {'sum': 140, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b01001011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2446,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 140, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011010; b = 8'b10001001; cin = 1'b1; // Expected: {'sum': 36, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011010; b = 8'b10001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2447,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 36, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b00101111; cin = 1'b0; // Expected: {'sum': 146, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b00101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2448,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 146, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b10111101; cin = 1'b1; // Expected: {'sum': 11, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b10111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2449,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 11, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011001; b = 8'b11000101; cin = 1'b0; // Expected: {'sum': 222, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011001; b = 8'b11000101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2450,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 222, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001111; b = 8'b10101110; cin = 1'b1; // Expected: {'sum': 254, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001111; b = 8'b10101110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2451,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 254, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b01010110; cin = 1'b1; // Expected: {'sum': 233, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b01010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2452,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 233, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b01111000; cin = 1'b0; // Expected: {'sum': 108, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b01111000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2453,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 108, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110100; b = 8'b10010000; cin = 1'b0; // Expected: {'sum': 4, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110100; b = 8'b10010000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2454,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b01000100; cin = 1'b1; // Expected: {'sum': 160, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b01000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2455,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 160, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b00011000; cin = 1'b0; // Expected: {'sum': 165, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b00011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2456,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 165, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b10100011; cin = 1'b0; // Expected: {'sum': 59, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b10100011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2457,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 59, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b10010111; cin = 1'b0; // Expected: {'sum': 170, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b10010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2458,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 170, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b01001011; cin = 1'b0; // Expected: {'sum': 214, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b01001011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2459,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 214, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b10001101; cin = 1'b0; // Expected: {'sum': 40, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b10001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2460,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 40, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b11010101; cin = 1'b1; // Expected: {'sum': 165, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b11010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2461,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 165, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b11101110; cin = 1'b0; // Expected: {'sum': 224, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b11101110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2462,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 224, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b10100101; cin = 1'b0; // Expected: {'sum': 158, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b10100101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2463,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 158, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010100; b = 8'b10110100; cin = 1'b0; // Expected: {'sum': 200, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010100; b = 8'b10110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2464,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 200, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b00101011; cin = 1'b1; // Expected: {'sum': 120, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b00101011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2465,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 120, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110000; b = 8'b00010000; cin = 1'b1; // Expected: {'sum': 65, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110000; b = 8'b00010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2466,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 65, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b11111110; cin = 1'b1; // Expected: {'sum': 53, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b11111110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2467,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 53, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b11100110; cin = 1'b1; // Expected: {'sum': 5, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b11100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2468,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 5, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011100; b = 8'b00010011; cin = 1'b0; // Expected: {'sum': 239, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011100; b = 8'b00010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2469,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 239, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b11100111; cin = 1'b1; // Expected: {'sum': 213, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b11100111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2470,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 213, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b10011000; cin = 1'b0; // Expected: {'sum': 138, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b10011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2471,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 138, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b01100110; cin = 1'b0; // Expected: {'sum': 188, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b01100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2472,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 188, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b00100010; cin = 1'b0; // Expected: {'sum': 178, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b00100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2473,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 178, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b11000101; cin = 1'b1; // Expected: {'sum': 69, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b11000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2474,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 69, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b10101111; cin = 1'b1; // Expected: {'sum': 59, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b10101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2475,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 59, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b01010011; cin = 1'b1; // Expected: {'sum': 35, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b01010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2476,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 35, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111111; b = 8'b10001110; cin = 1'b0; // Expected: {'sum': 205, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111111; b = 8'b10001110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2477,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 205, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110011; b = 8'b00011100; cin = 1'b1; // Expected: {'sum': 208, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110011; b = 8'b00011100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2478,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 208, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001100; b = 8'b10001101; cin = 1'b0; // Expected: {'sum': 25, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001100; b = 8'b10001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2479,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 25, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001101; b = 8'b10010011; cin = 1'b1; // Expected: {'sum': 97, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001101; b = 8'b10010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2480,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 97, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b01111100; cin = 1'b1; // Expected: {'sum': 142, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b01111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2481,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 142, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000110; b = 8'b10111110; cin = 1'b0; // Expected: {'sum': 196, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000110; b = 8'b10111110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2482,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 196, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b00111111; cin = 1'b0; // Expected: {'sum': 187, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b00111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2483,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 187, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b00100011; cin = 1'b0; // Expected: {'sum': 86, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b00100011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2484,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 86, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b10011111; cin = 1'b0; // Expected: {'sum': 158, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b10011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2485,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 158, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101111; b = 8'b10000111; cin = 1'b1; // Expected: {'sum': 247, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101111; b = 8'b10000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2486,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 247, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100001; b = 8'b00010010; cin = 1'b0; // Expected: {'sum': 51, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100001; b = 8'b00010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2487,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 51, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b10111001; cin = 1'b0; // Expected: {'sum': 209, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b10111001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2488,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 209, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b00110111; cin = 1'b1; // Expected: {'sum': 58, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b00110111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2489,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 58, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011010; b = 8'b10111110; cin = 1'b0; // Expected: {'sum': 88, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011010; b = 8'b10111110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2490,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 88, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110100; b = 8'b10111001; cin = 1'b0; // Expected: {'sum': 45, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110100; b = 8'b10111001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2491,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 45, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b00010110; cin = 1'b1; // Expected: {'sum': 248, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b00010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2492,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 248, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b11001110; cin = 1'b1; // Expected: {'sum': 97, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b11001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2493,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 97, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b01011011; cin = 1'b0; // Expected: {'sum': 171, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b01011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2494,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 171, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b01010011; cin = 1'b0; // Expected: {'sum': 163, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b01010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2495,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 163, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010100; b = 8'b10010110; cin = 1'b1; // Expected: {'sum': 107, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010100; b = 8'b10010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2496,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 107, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b00111100; cin = 1'b0; // Expected: {'sum': 190, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b00111100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2497,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 190, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b00011111; cin = 1'b0; // Expected: {'sum': 22, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b00011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2498,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 22, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b01101101; cin = 1'b1; // Expected: {'sum': 196, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b01101101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2499,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 196, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b01111111; cin = 1'b0; // Expected: {'sum': 161, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b01111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2500,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 161, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b00000001; cin = 1'b0; // Expected: {'sum': 208, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b00000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2501,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 208, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b10111000; cin = 1'b1; // Expected: {'sum': 49, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b10111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2502,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 49, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b10011010; cin = 1'b1; // Expected: {'sum': 55, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b10011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2503,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 55, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101110; b = 8'b00001000; cin = 1'b0; // Expected: {'sum': 54, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101110; b = 8'b00001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2504,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 54, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b00011000; cin = 1'b1; // Expected: {'sum': 70, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b00011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2505,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 70, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b11111111; cin = 1'b0; // Expected: {'sum': 125, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b11111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2506,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 125, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000111; b = 8'b11100010; cin = 1'b1; // Expected: {'sum': 170, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000111; b = 8'b11100010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2507,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 170, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b00111111; cin = 1'b1; // Expected: {'sum': 141, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b00111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2508,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 141, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100000; b = 8'b11011001; cin = 1'b0; // Expected: {'sum': 57, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100000; b = 8'b11011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2509,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 57, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010011; b = 8'b11011001; cin = 1'b0; // Expected: {'sum': 172, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010011; b = 8'b11011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2510,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 172, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b10111011; cin = 1'b0; // Expected: {'sum': 116, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b10111011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2511,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 116, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000110; b = 8'b10001100; cin = 1'b1; // Expected: {'sum': 147, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000110; b = 8'b10001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2512,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 147, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b11010100; cin = 1'b1; // Expected: {'sum': 100, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b11010100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2513,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 100, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b01010010; cin = 1'b0; // Expected: {'sum': 113, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b01010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2514,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 113, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b10001100; cin = 1'b1; // Expected: {'sum': 176, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b10001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2515,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 176, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100001; b = 8'b11111000; cin = 1'b0; // Expected: {'sum': 25, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100001; b = 8'b11111000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2516,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 25, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b11010011; cin = 1'b1; // Expected: {'sum': 132, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b11010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2517,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 132, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101000; b = 8'b10111111; cin = 1'b0; // Expected: {'sum': 231, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101000; b = 8'b10111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2518,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 231, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011000; b = 8'b00011011; cin = 1'b0; // Expected: {'sum': 115, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011000; b = 8'b00011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2519,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 115, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b01000010; cin = 1'b0; // Expected: {'sum': 85, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b01000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2520,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 85, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b01010110; cin = 1'b1; // Expected: {'sum': 38, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b01010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2521,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 38, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b00101010; cin = 1'b0; // Expected: {'sum': 92, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b00101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2522,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 92, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100010; b = 8'b00001000; cin = 1'b1; // Expected: {'sum': 235, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100010; b = 8'b00001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2523,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 235, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b11001100; cin = 1'b1; // Expected: {'sum': 42, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b11001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2524,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 42, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101010; b = 8'b00101111; cin = 1'b1; // Expected: {'sum': 26, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101010; b = 8'b00101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2525,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 26, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000001; b = 8'b10110101; cin = 1'b0; // Expected: {'sum': 118, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000001; b = 8'b10110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2526,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 118, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b10101010; cin = 1'b1; // Expected: {'sum': 84, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b10101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2527,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 84, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b00011011; cin = 1'b0; // Expected: {'sum': 13, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b00011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2528,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 13, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b11011001; cin = 1'b1; // Expected: {'sum': 208, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b11011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2529,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 208, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b01011010; cin = 1'b0; // Expected: {'sum': 212, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b01011010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2530,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 212, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b01010111; cin = 1'b1; // Expected: {'sum': 251, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b01010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2531,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 251, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b11011000; cin = 1'b0; // Expected: {'sum': 247, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b11011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2532,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 247, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001011; b = 8'b01110100; cin = 1'b1; // Expected: {'sum': 128, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001011; b = 8'b01110100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2533,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 128, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b10101001; cin = 1'b0; // Expected: {'sum': 44, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b10101001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2534,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 44, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100000; b = 8'b10010111; cin = 1'b0; // Expected: {'sum': 247, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100000; b = 8'b10010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2535,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 247, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010110; b = 8'b01001100; cin = 1'b0; // Expected: {'sum': 34, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010110; b = 8'b01001100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2536,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 34, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001110; b = 8'b11011011; cin = 1'b0; // Expected: {'sum': 233, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001110; b = 8'b11011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2537,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 233, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b00011101; cin = 1'b0; // Expected: {'sum': 24, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b00011101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2538,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 24, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100000; b = 8'b11010111; cin = 1'b0; // Expected: {'sum': 55, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100000; b = 8'b11010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2539,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 55, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001011; b = 8'b11111111; cin = 1'b1; // Expected: {'sum': 75, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001011; b = 8'b11111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2540,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 75, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011111; b = 8'b11101110; cin = 1'b0; // Expected: {'sum': 77, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011111; b = 8'b11101110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2541,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 77, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111010; b = 8'b11100101; cin = 1'b1; // Expected: {'sum': 224, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111010; b = 8'b11100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2542,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 224, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b11111101; cin = 1'b0; // Expected: {'sum': 143, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b11111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2543,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 143, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b00101100; cin = 1'b0; // Expected: {'sum': 39, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b00101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2544,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 39, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b10100010; cin = 1'b1; // Expected: {'sum': 173, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b10100010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2545,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 173, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b11011001; cin = 1'b1; // Expected: {'sum': 68, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b11011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2546,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 68, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010011; b = 8'b00111101; cin = 1'b1; // Expected: {'sum': 17, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010011; b = 8'b00111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2547,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 17, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b01010100; cin = 1'b0; // Expected: {'sum': 92, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b01010100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2548,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 92, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000111; b = 8'b00011011; cin = 1'b1; // Expected: {'sum': 163, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000111; b = 8'b00011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2549,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 163, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b01110111; cin = 1'b0; // Expected: {'sum': 241, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b01110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2550,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 241, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b10010010; cin = 1'b1; // Expected: {'sum': 212, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b10010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2551,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 212, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000100; b = 8'b11000111; cin = 1'b1; // Expected: {'sum': 204, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000100; b = 8'b11000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2552,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 204, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101001; b = 8'b01111001; cin = 1'b1; // Expected: {'sum': 227, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101001; b = 8'b01111001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2553,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 227, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b11100111; cin = 1'b1; // Expected: {'sum': 68, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b11100111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2554,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 68, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b01101000; cin = 1'b1; // Expected: {'sum': 84, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b01101000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2555,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 84, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000011; b = 8'b10111101; cin = 1'b1; // Expected: {'sum': 129, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000011; b = 8'b10111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2556,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 129, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b10101011; cin = 1'b0; // Expected: {'sum': 140, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b10101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2557,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 140, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101100; b = 8'b10101100; cin = 1'b0; // Expected: {'sum': 152, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101100; b = 8'b10101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2558,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 152, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b11111100; cin = 1'b1; // Expected: {'sum': 49, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b11111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2559,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 49, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010111; b = 8'b10011100; cin = 1'b1; // Expected: {'sum': 244, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010111; b = 8'b10011100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2560,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 244, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011010; b = 8'b11010010; cin = 1'b1; // Expected: {'sum': 45, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011010; b = 8'b11010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2561,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 45, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111111; b = 8'b10000001; cin = 1'b1; // Expected: {'sum': 193, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111111; b = 8'b10000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2562,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 193, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b00110010; cin = 1'b0; // Expected: {'sum': 148, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b00110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2563,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 148, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b01110001; cin = 1'b0; // Expected: {'sum': 158, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b01110001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2564,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 158, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b10101111; cin = 1'b1; // Expected: {'sum': 241, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b10101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2565,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 241, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b00001100; cin = 1'b1; // Expected: {'sum': 110, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b00001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2566,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 110, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001101; b = 8'b00100111; cin = 1'b0; // Expected: {'sum': 244, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001101; b = 8'b00100111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2567,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 244, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b01101111; cin = 1'b1; // Expected: {'sum': 21, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b01101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2568,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 21, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110001; b = 8'b01111100; cin = 1'b0; // Expected: {'sum': 173, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110001; b = 8'b01111100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2569,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 173, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111111; b = 8'b01011101; cin = 1'b0; // Expected: {'sum': 156, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111111; b = 8'b01011101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2570,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 156, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001010; b = 8'b01100000; cin = 1'b1; // Expected: {'sum': 235, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001010; b = 8'b01100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2571,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 235, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b01011100; cin = 1'b0; // Expected: {'sum': 71, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b01011100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2572,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 71, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001010; b = 8'b00100100; cin = 1'b1; // Expected: {'sum': 175, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001010; b = 8'b00100100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2573,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 175, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010000; b = 8'b01100101; cin = 1'b1; // Expected: {'sum': 118, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010000; b = 8'b01100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2574,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 118, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b00010011; cin = 1'b0; // Expected: {'sum': 36, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b00010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2575,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 36, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b11010011; cin = 1'b0; // Expected: {'sum': 75, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b11010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2576,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 75, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011001; b = 8'b00110110; cin = 1'b1; // Expected: {'sum': 208, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011001; b = 8'b00110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2577,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 208, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b10010100; cin = 1'b1; // Expected: {'sum': 39, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b10010100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2578,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 39, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b10101011; cin = 1'b1; // Expected: {'sum': 141, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b10101011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2579,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 141, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b00011001; cin = 1'b1; // Expected: {'sum': 187, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b00011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2580,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 187, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b00001011; cin = 1'b0; // Expected: {'sum': 11, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b00001011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2581,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 11, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010010; b = 8'b01000101; cin = 1'b1; // Expected: {'sum': 152, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010010; b = 8'b01000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2582,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 152, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b10011111; cin = 1'b1; // Expected: {'sum': 123, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b10011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2583,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 123, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b11010101; cin = 1'b0; // Expected: {'sum': 82, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b11010101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2584,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 82, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b00101000; cin = 1'b0; // Expected: {'sum': 77, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b00101000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2585,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 77, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b00001100; cin = 1'b1; // Expected: {'sum': 199, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b00001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2586,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 199, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b01000100; cin = 1'b1; // Expected: {'sum': 121, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b01000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2587,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 121, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100111; b = 8'b01010101; cin = 1'b1; // Expected: {'sum': 253, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100111; b = 8'b01010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2588,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 253, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001011; b = 8'b00011000; cin = 1'b0; // Expected: {'sum': 35, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001011; b = 8'b00011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2589,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 35, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b10101011; cin = 1'b0; // Expected: {'sum': 251, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b10101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2590,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 251, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010000; b = 8'b01111110; cin = 1'b0; // Expected: {'sum': 142, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010000; b = 8'b01111110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2591,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 142, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b00110111; cin = 1'b1; // Expected: {'sum': 64, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b00110111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2592,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 64, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b10101001; cin = 1'b0; // Expected: {'sum': 58, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b10101001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2593,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 58, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b10011000; cin = 1'b0; // Expected: {'sum': 218, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b10011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2594,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 218, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010110; b = 8'b01001101; cin = 1'b0; // Expected: {'sum': 35, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010110; b = 8'b01001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2595,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 35, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111101; b = 8'b10010001; cin = 1'b0; // Expected: {'sum': 206, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111101; b = 8'b10010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2596,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 206, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101110; b = 8'b10000010; cin = 1'b1; // Expected: {'sum': 177, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101110; b = 8'b10000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2597,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 177, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b00011100; cin = 1'b1; // Expected: {'sum': 198, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b00011100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2598,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 198, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b11111011; cin = 1'b0; // Expected: {'sum': 110, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b11111011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2599,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 110, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b11011010; cin = 1'b0; // Expected: {'sum': 88, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b11011010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2600,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 88, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b11101111; cin = 1'b1; // Expected: {'sum': 7, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b11101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2601,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001001; b = 8'b11111000; cin = 1'b0; // Expected: {'sum': 65, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001001; b = 8'b11111000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2602,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 65, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b10100000; cin = 1'b1; // Expected: {'sum': 150, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b10100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2603,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 150, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b11110110; cin = 1'b1; // Expected: {'sum': 235, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b11110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2604,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 235, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b00101100; cin = 1'b1; // Expected: {'sum': 175, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b00101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2605,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 175, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b10000010; cin = 1'b1; // Expected: {'sum': 148, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b10000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2606,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 148, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b10111000; cin = 1'b1; // Expected: {'sum': 170, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b10111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2607,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 170, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000111; b = 8'b01100010; cin = 1'b0; // Expected: {'sum': 41, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000111; b = 8'b01100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2608,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 41, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010010; b = 8'b11001000; cin = 1'b0; // Expected: {'sum': 26, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010010; b = 8'b11001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2609,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 26, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b00011011; cin = 1'b1; // Expected: {'sum': 234, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b00011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2610,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 234, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b01000011; cin = 1'b0; // Expected: {'sum': 230, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b01000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2611,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 230, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110110; b = 8'b11010110; cin = 1'b0; // Expected: {'sum': 76, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110110; b = 8'b11010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2612,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 76, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111110; b = 8'b00111101; cin = 1'b1; // Expected: {'sum': 124, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111110; b = 8'b00111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2613,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 124, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b11101100; cin = 1'b1; // Expected: {'sum': 89, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b11101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2614,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 89, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b00101100; cin = 1'b0; // Expected: {'sum': 189, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b00101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2615,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 189, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b11011001; cin = 1'b0; // Expected: {'sum': 139, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b11011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2616,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 139, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111000; b = 8'b11001000; cin = 1'b0; // Expected: {'sum': 0, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111000; b = 8'b11001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2617,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b00100011; cin = 1'b0; // Expected: {'sum': 20, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b00100011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2618,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 20, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b00001010; cin = 1'b0; // Expected: {'sum': 185, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b00001010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2619,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 185, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111101; b = 8'b11100000; cin = 1'b1; // Expected: {'sum': 30, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111101; b = 8'b11100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2620,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 30, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b11011110; cin = 1'b1; // Expected: {'sum': 144, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b11011110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2621,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 144, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b11010011; cin = 1'b0; // Expected: {'sum': 131, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b11010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2622,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 131, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010010; b = 8'b11100101; cin = 1'b0; // Expected: {'sum': 247, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010010; b = 8'b11100101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2623,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 247, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b11101001; cin = 1'b1; // Expected: {'sum': 43, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b11101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2624,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 43, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b10111111; cin = 1'b0; // Expected: {'sum': 29, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b10111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2625,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 29, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b01001101; cin = 1'b0; // Expected: {'sum': 183, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b01001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2626,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 183, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111010; b = 8'b11110000; cin = 1'b1; // Expected: {'sum': 235, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111010; b = 8'b11110000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2627,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 235, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b11000001; cin = 1'b1; // Expected: {'sum': 101, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b11000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2628,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 101, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b10001000; cin = 1'b0; // Expected: {'sum': 0, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b10001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2629,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b00101111; cin = 1'b0; // Expected: {'sum': 33, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b00101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2630,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 33, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110101; b = 8'b11111111; cin = 1'b1; // Expected: {'sum': 181, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110101; b = 8'b11111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2631,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 181, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b10100110; cin = 1'b1; // Expected: {'sum': 202, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b10100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2632,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 202, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b01010001; cin = 1'b1; // Expected: {'sum': 242, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b01010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2633,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 242, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b00111101; cin = 1'b1; // Expected: {'sum': 223, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b00111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2634,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 223, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b11101001; cin = 1'b0; // Expected: {'sum': 171, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b11101001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2635,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 171, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b01100110; cin = 1'b1; // Expected: {'sum': 60, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b01100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2636,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 60, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b11000010; cin = 1'b1; // Expected: {'sum': 245, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b11000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2637,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 245, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011010; b = 8'b10001101; cin = 1'b1; // Expected: {'sum': 104, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011010; b = 8'b10001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2638,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 104, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b10011000; cin = 1'b0; // Expected: {'sum': 33, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b10011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2639,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 33, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b10111001; cin = 1'b0; // Expected: {'sum': 29, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b10111001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2640,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 29, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b01001100; cin = 1'b1; // Expected: {'sum': 66, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b01001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2641,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 66, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b01000100; cin = 1'b0; // Expected: {'sum': 68, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b01000100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2642,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 68, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b00000010; cin = 1'b1; // Expected: {'sum': 122, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b00000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2643,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 122, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b01001011; cin = 1'b0; // Expected: {'sum': 104, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b01001011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2644,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 104, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b10100100; cin = 1'b0; // Expected: {'sum': 173, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b10100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2645,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 173, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b10000001; cin = 1'b0; // Expected: {'sum': 194, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b10000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2646,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 194, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001000; b = 8'b11010011; cin = 1'b1; // Expected: {'sum': 28, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001000; b = 8'b11010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2647,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 28, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b10111001; cin = 1'b0; // Expected: {'sum': 9, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b10111001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2648,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 9, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b00101011; cin = 1'b0; // Expected: {'sum': 30, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b00101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2649,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 30, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b11010001; cin = 1'b1; // Expected: {'sum': 209, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b11010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2650,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 209, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100110; b = 8'b10110010; cin = 1'b1; // Expected: {'sum': 153, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100110; b = 8'b10110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2651,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 153, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b00000101; cin = 1'b0; // Expected: {'sum': 42, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b00000101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2652,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 42, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b10101011; cin = 1'b0; // Expected: {'sum': 125, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b10101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2653,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 125, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100111; b = 8'b10111101; cin = 1'b1; // Expected: {'sum': 37, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100111; b = 8'b10111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2654,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 37, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b01011000; cin = 1'b1; // Expected: {'sum': 27, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b01011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2655,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 27, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100100; b = 8'b11011100; cin = 1'b1; // Expected: {'sum': 129, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100100; b = 8'b11011100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2656,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 129, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001100; b = 8'b11000100; cin = 1'b0; // Expected: {'sum': 80, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001100; b = 8'b11000100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2657,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 80, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b00111000; cin = 1'b0; // Expected: {'sum': 15, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b00111000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2658,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b11000011; cin = 1'b0; // Expected: {'sum': 75, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b11000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2659,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 75, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b11000110; cin = 1'b0; // Expected: {'sum': 232, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b11000110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2660,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 232, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b11100001; cin = 1'b1; // Expected: {'sum': 211, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b11100001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2661,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 211, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b00010000; cin = 1'b1; // Expected: {'sum': 183, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b00010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2662,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 183, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b00001110; cin = 1'b1; // Expected: {'sum': 1, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b00001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2663,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b11100111; cin = 1'b0; // Expected: {'sum': 33, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b11100111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2664,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 33, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b01100011; cin = 1'b1; // Expected: {'sum': 165, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b01100011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2665,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 165, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b00111010; cin = 1'b1; // Expected: {'sum': 43, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b00111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2666,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 43, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b11111001; cin = 1'b1; // Expected: {'sum': 20, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b11111001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2667,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 20, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b01101011; cin = 1'b0; // Expected: {'sum': 57, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b01101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2668,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 57, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011101; b = 8'b00000101; cin = 1'b1; // Expected: {'sum': 163, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011101; b = 8'b00000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2669,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 163, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100000; b = 8'b01010110; cin = 1'b0; // Expected: {'sum': 54, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100000; b = 8'b01010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2670,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 54, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b01100000; cin = 1'b0; // Expected: {'sum': 161, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b01100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2671,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 161, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b10111001; cin = 1'b1; // Expected: {'sum': 6, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b10111001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2672,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b10001100; cin = 1'b1; // Expected: {'sum': 201, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b10001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2673,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 201, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b11010110; cin = 1'b1; // Expected: {'sum': 194, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b11010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2674,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 194, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b11100100; cin = 1'b1; // Expected: {'sum': 14, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b11100100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2675,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110101; b = 8'b11111001; cin = 1'b1; // Expected: {'sum': 175, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110101; b = 8'b11111001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2676,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 175, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b01101010; cin = 1'b1; // Expected: {'sum': 157, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b01101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2677,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 157, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b01000000; cin = 1'b1; // Expected: {'sum': 16, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b01000000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2678,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 16, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b11110101; cin = 1'b0; // Expected: {'sum': 238, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b11110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2679,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 238, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b11011001; cin = 1'b0; // Expected: {'sum': 222, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b11011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2680,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 222, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b01000001; cin = 1'b0; // Expected: {'sum': 215, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b01000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2681,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 215, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b00001000; cin = 1'b0; // Expected: {'sum': 152, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b00001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2682,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 152, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b11010001; cin = 1'b0; // Expected: {'sum': 33, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b11010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2683,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 33, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000011; b = 8'b01011101; cin = 1'b0; // Expected: {'sum': 32, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000011; b = 8'b01011101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2684,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 32, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b10011000; cin = 1'b1; // Expected: {'sum': 153, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b10011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2685,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 153, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b01111010; cin = 1'b1; // Expected: {'sum': 175, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b01111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2686,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 175, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100000; b = 8'b10011001; cin = 1'b0; // Expected: {'sum': 185, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100000; b = 8'b10011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2687,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 185, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b00010100; cin = 1'b1; // Expected: {'sum': 51, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b00010100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2688,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 51, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b01011010; cin = 1'b1; // Expected: {'sum': 80, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b01011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2689,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 80, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b10101011; cin = 1'b1; // Expected: {'sum': 161, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b10101011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2690,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 161, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b11110110; cin = 1'b0; // Expected: {'sum': 206, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b11110110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2691,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 206, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b11000100; cin = 1'b1; // Expected: {'sum': 204, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b11000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2692,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 204, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b00001011; cin = 1'b1; // Expected: {'sum': 92, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b00001011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2693,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 92, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b10101001; cin = 1'b1; // Expected: {'sum': 35, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b10101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2694,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 35, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b11010110; cin = 1'b1; // Expected: {'sum': 210, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b11010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2695,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 210, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b01010111; cin = 1'b0; // Expected: {'sum': 46, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b01010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2696,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 46, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000001; b = 8'b10110100; cin = 1'b1; // Expected: {'sum': 118, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000001; b = 8'b10110100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2697,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 118, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b01100110; cin = 1'b0; // Expected: {'sum': 22, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b01100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2698,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 22, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b01101011; cin = 1'b1; // Expected: {'sum': 225, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b01101011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2699,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 225, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b11110010; cin = 1'b0; // Expected: {'sum': 142, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b11110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2700,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 142, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100111; b = 8'b10001011; cin = 1'b0; // Expected: {'sum': 50, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100111; b = 8'b10001011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2701,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 50, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011000; b = 8'b10001110; cin = 1'b0; // Expected: {'sum': 230, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011000; b = 8'b10001110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2702,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 230, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101001; b = 8'b00100111; cin = 1'b1; // Expected: {'sum': 17, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101001; b = 8'b00100111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2703,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 17, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b10101111; cin = 1'b0; // Expected: {'sum': 46, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b10101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2704,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 46, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b10000000; cin = 1'b0; // Expected: {'sum': 118, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b10000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2705,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 118, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b00111111; cin = 1'b1; // Expected: {'sum': 205, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b00111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2706,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 205, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001101; b = 8'b00001110; cin = 1'b1; // Expected: {'sum': 220, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001101; b = 8'b00001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2707,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 220, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b11101110; cin = 1'b1; // Expected: {'sum': 185, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b11101110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2708,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 185, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001110; b = 8'b10000000; cin = 1'b1; // Expected: {'sum': 207, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001110; b = 8'b10000000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2709,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 207, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b01000001; cin = 1'b1; // Expected: {'sum': 27, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b01000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2710,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 27, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101111; b = 8'b01110110; cin = 1'b1; // Expected: {'sum': 166, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101111; b = 8'b01110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2711,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 166, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010011; b = 8'b10100011; cin = 1'b0; // Expected: {'sum': 246, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010011; b = 8'b10100011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2712,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 246, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b01001001; cin = 1'b0; // Expected: {'sum': 199, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b01001001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2713,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 199, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000110; b = 8'b01010111; cin = 1'b0; // Expected: {'sum': 157, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000110; b = 8'b01010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2714,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 157, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101111; b = 8'b11001010; cin = 1'b1; // Expected: {'sum': 250, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101111; b = 8'b11001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2715,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 250, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b10100111; cin = 1'b0; // Expected: {'sum': 227, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b10100111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2716,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 227, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011011; b = 8'b01001010; cin = 1'b0; // Expected: {'sum': 101, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011011; b = 8'b01001010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2717,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 101, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b11010101; cin = 1'b0; // Expected: {'sum': 65, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b11010101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2718,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 65, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b10100010; cin = 1'b0; // Expected: {'sum': 167, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b10100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2719,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 167, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101111; b = 8'b00010011; cin = 1'b0; // Expected: {'sum': 66, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101111; b = 8'b00010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2720,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 66, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b01110011; cin = 1'b1; // Expected: {'sum': 52, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b01110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2721,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 52, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b10111101; cin = 1'b0; // Expected: {'sum': 185, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b10111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2722,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 185, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010100; b = 8'b01101111; cin = 1'b1; // Expected: {'sum': 132, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010100; b = 8'b01101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2723,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 132, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b11100101; cin = 1'b1; // Expected: {'sum': 202, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b11100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2724,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 202, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111011; b = 8'b00000101; cin = 1'b0; // Expected: {'sum': 128, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111011; b = 8'b00000101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2725,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 128, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011111; b = 8'b00001111; cin = 1'b1; // Expected: {'sum': 111, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011111; b = 8'b00001111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2726,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 111, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b00110000; cin = 1'b0; // Expected: {'sum': 237, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b00110000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2727,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 237, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b10100001; cin = 1'b1; // Expected: {'sum': 185, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b10100001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2728,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 185, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b11101010; cin = 1'b1; // Expected: {'sum': 47, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b11101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2729,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 47, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b11010001; cin = 1'b0; // Expected: {'sum': 94, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b11010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2730,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 94, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000000; b = 8'b01001001; cin = 1'b0; // Expected: {'sum': 201, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000000; b = 8'b01001001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2731,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 201, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000110; b = 8'b01001011; cin = 1'b1; // Expected: {'sum': 146, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000110; b = 8'b01001011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2732,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 146, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100110; b = 8'b10001111; cin = 1'b0; // Expected: {'sum': 181, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100110; b = 8'b10001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2733,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 181, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b01100101; cin = 1'b0; // Expected: {'sum': 68, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b01100101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2734,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 68, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b10010001; cin = 1'b0; // Expected: {'sum': 195, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b10010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2735,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 195, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b01101000; cin = 1'b1; // Expected: {'sum': 115, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b01101000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2736,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 115, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001011; b = 8'b01010111; cin = 1'b1; // Expected: {'sum': 35, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001011; b = 8'b01010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2737,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 35, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b00000001; cin = 1'b0; // Expected: {'sum': 162, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b00000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2738,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 162, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b01110010; cin = 1'b1; // Expected: {'sum': 237, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b01110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2739,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 237, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b01011111; cin = 1'b1; // Expected: {'sum': 83, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b01011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2740,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 83, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b01110011; cin = 1'b0; // Expected: {'sum': 156, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b01110011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2741,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 156, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001100; b = 8'b00110101; cin = 1'b0; // Expected: {'sum': 193, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001100; b = 8'b00110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2742,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 193, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b11010000; cin = 1'b0; // Expected: {'sum': 225, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b11010000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2743,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 225, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000111; b = 8'b11001110; cin = 1'b0; // Expected: {'sum': 149, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000111; b = 8'b11001110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2744,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 149, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100111; b = 8'b00111111; cin = 1'b1; // Expected: {'sum': 39, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100111; b = 8'b00111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2745,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 39, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100110; b = 8'b01111100; cin = 1'b1; // Expected: {'sum': 227, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100110; b = 8'b01111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2746,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 227, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101010; b = 8'b00010010; cin = 1'b0; // Expected: {'sum': 252, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101010; b = 8'b00010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2747,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 252, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001111; b = 8'b10000111; cin = 1'b1; // Expected: {'sum': 151, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001111; b = 8'b10000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2748,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 151, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b11111010; cin = 1'b0; // Expected: {'sum': 209, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b11111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2749,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 209, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b11010001; cin = 1'b0; // Expected: {'sum': 52, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b11010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2750,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 52, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b10010101; cin = 1'b1; // Expected: {'sum': 16, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b10010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2751,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 16, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b01100110; cin = 1'b0; // Expected: {'sum': 224, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b01100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2752,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 224, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101101; b = 8'b10010011; cin = 1'b1; // Expected: {'sum': 65, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101101; b = 8'b10010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2753,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 65, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b01111100; cin = 1'b1; // Expected: {'sum': 252, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b01111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2754,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 252, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b11011111; cin = 1'b1; // Expected: {'sum': 87, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b11011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2755,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 87, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b00111100; cin = 1'b1; // Expected: {'sum': 21, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b00111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2756,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 21, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011011; b = 8'b00011000; cin = 1'b1; // Expected: {'sum': 52, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011011; b = 8'b00011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2757,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 52, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110001; b = 8'b11000010; cin = 1'b1; // Expected: {'sum': 244, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110001; b = 8'b11000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2758,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 244, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b01110101; cin = 1'b0; // Expected: {'sum': 182, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b01110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2759,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 182, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b11101010; cin = 1'b1; // Expected: {'sum': 46, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b11101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2760,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 46, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b00011110; cin = 1'b0; // Expected: {'sum': 53, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b00011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2761,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 53, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100010; b = 8'b01010111; cin = 1'b0; // Expected: {'sum': 57, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100010; b = 8'b01010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2762,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 57, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b11100011; cin = 1'b0; // Expected: {'sum': 92, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b11100011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2763,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 92, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000111; b = 8'b00000001; cin = 1'b1; // Expected: {'sum': 201, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000111; b = 8'b00000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2764,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 201, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b11011101; cin = 1'b1; // Expected: {'sum': 122, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b11011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2765,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 122, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000101; b = 8'b10000110; cin = 1'b1; // Expected: {'sum': 12, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000101; b = 8'b10000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2766,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b00111111; cin = 1'b1; // Expected: {'sum': 198, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b00111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2767,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 198, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b10101101; cin = 1'b1; // Expected: {'sum': 167, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b10101101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2768,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 167, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b00111011; cin = 1'b1; // Expected: {'sum': 91, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b00111011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2769,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 91, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b00011011; cin = 1'b0; // Expected: {'sum': 16, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b00011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2770,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 16, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000001; b = 8'b10001001; cin = 1'b1; // Expected: {'sum': 75, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000001; b = 8'b10001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2771,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 75, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b01000100; cin = 1'b0; // Expected: {'sum': 134, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b01000100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2772,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 134, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b00011101; cin = 1'b1; // Expected: {'sum': 101, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b00011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2773,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 101, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b11001000; cin = 1'b1; // Expected: {'sum': 194, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b11001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2774,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 194, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011001; b = 8'b11011000; cin = 1'b0; // Expected: {'sum': 241, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011001; b = 8'b11011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2775,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 241, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b01100110; cin = 1'b0; // Expected: {'sum': 239, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b01100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2776,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 239, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b00110110; cin = 1'b1; // Expected: {'sum': 90, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b00110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2777,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 90, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b01101111; cin = 1'b0; // Expected: {'sum': 32, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b01101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2778,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 32, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001011; b = 8'b11000010; cin = 1'b1; // Expected: {'sum': 14, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001011; b = 8'b11000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2779,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101010; b = 8'b10000100; cin = 1'b1; // Expected: {'sum': 47, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101010; b = 8'b10000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2780,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 47, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011110; b = 8'b00011101; cin = 1'b0; // Expected: {'sum': 251, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011110; b = 8'b00011101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2781,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 251, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101111; b = 8'b00011111; cin = 1'b0; // Expected: {'sum': 142, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101111; b = 8'b00011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2782,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 142, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b10100000; cin = 1'b1; // Expected: {'sum': 219, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b10100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2783,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 219, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b10000011; cin = 1'b0; // Expected: {'sum': 166, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b10000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2784,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 166, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b11011010; cin = 1'b0; // Expected: {'sum': 205, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b11011010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2785,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 205, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b11011100; cin = 1'b1; // Expected: {'sum': 222, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b11011100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2786,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 222, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110110; b = 8'b10010111; cin = 1'b1; // Expected: {'sum': 14, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110110; b = 8'b10010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2787,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b11001000; cin = 1'b0; // Expected: {'sum': 173, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b11001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2788,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 173, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b10010111; cin = 1'b1; // Expected: {'sum': 3, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b10010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2789,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010011; b = 8'b11011000; cin = 1'b1; // Expected: {'sum': 108, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010011; b = 8'b11011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2790,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 108, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b11000011; cin = 1'b0; // Expected: {'sum': 193, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b11000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2791,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 193, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b10111011; cin = 1'b0; // Expected: {'sum': 150, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b10111011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2792,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 150, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b00111110; cin = 1'b1; // Expected: {'sum': 39, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b00111110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2793,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 39, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b11110101; cin = 1'b1; // Expected: {'sum': 186, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b11110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2794,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 186, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011011; b = 8'b10000110; cin = 1'b1; // Expected: {'sum': 162, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011011; b = 8'b10000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2795,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 162, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b01100110; cin = 1'b1; // Expected: {'sum': 189, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b01100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2796,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 189, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b01100111; cin = 1'b1; // Expected: {'sum': 50, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b01100111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2797,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 50, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b00100001; cin = 1'b0; // Expected: {'sum': 250, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b00100001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2798,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 250, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b10000101; cin = 1'b1; // Expected: {'sum': 220, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b10000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2799,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 220, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b01101100; cin = 1'b0; // Expected: {'sum': 232, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b01101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2800,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 232, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b10001110; cin = 1'b1; // Expected: {'sum': 132, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b10001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2801,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 132, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000100; b = 8'b10100101; cin = 1'b1; // Expected: {'sum': 170, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000100; b = 8'b10100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2802,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 170, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b00101000; cin = 1'b1; // Expected: {'sum': 192, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b00101000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2803,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 192, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b11110100; cin = 1'b1; // Expected: {'sum': 197, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b11110100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2804,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 197, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b11001101; cin = 1'b1; // Expected: {'sum': 47, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b11001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2805,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 47, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b00001100; cin = 1'b0; // Expected: {'sum': 14, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b00001100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2806,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010011; b = 8'b00111100; cin = 1'b0; // Expected: {'sum': 207, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010011; b = 8'b00111100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2807,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 207, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001000; b = 8'b01110001; cin = 1'b1; // Expected: {'sum': 58, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001000; b = 8'b01110001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2808,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 58, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b10011110; cin = 1'b0; // Expected: {'sum': 223, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b10011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2809,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 223, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b11110110; cin = 1'b1; // Expected: {'sum': 84, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b11110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2810,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 84, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100111; b = 8'b11100111; cin = 1'b1; // Expected: {'sum': 143, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100111; b = 8'b11100111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2811,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 143, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101010; b = 8'b00100110; cin = 1'b1; // Expected: {'sum': 209, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101010; b = 8'b00100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2812,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 209, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b11100000; cin = 1'b0; // Expected: {'sum': 92, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b11100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2813,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 92, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b11101001; cin = 1'b0; // Expected: {'sum': 145, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b11101001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2814,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 145, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011111; b = 8'b11000000; cin = 1'b1; // Expected: {'sum': 32, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011111; b = 8'b11000000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2815,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 32, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111000; b = 8'b10001101; cin = 1'b1; // Expected: {'sum': 198, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111000; b = 8'b10001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2816,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 198, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b10010110; cin = 1'b0; // Expected: {'sum': 45, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b10010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2817,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 45, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b01010010; cin = 1'b1; // Expected: {'sum': 182, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b01010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2818,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 182, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001000; b = 8'b01101111; cin = 1'b1; // Expected: {'sum': 184, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001000; b = 8'b01101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2819,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 184, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b11001101; cin = 1'b1; // Expected: {'sum': 16, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b11001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2820,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 16, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b10010001; cin = 1'b1; // Expected: {'sum': 125, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b10010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2821,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 125, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001011; b = 8'b01001101; cin = 1'b1; // Expected: {'sum': 25, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001011; b = 8'b01001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2822,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 25, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010100; b = 8'b10001011; cin = 1'b0; // Expected: {'sum': 223, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010100; b = 8'b10001011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2823,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 223, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b10100010; cin = 1'b0; // Expected: {'sum': 233, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b10100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2824,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 233, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000000; b = 8'b10111000; cin = 1'b0; // Expected: {'sum': 56, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000000; b = 8'b10111000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2825,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 56, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b01111110; cin = 1'b1; // Expected: {'sum': 86, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b01111110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2826,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 86, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b11100101; cin = 1'b0; // Expected: {'sum': 44, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b11100101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2827,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 44, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b01010100; cin = 1'b1; // Expected: {'sum': 166, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b01010100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2828,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 166, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b00001101; cin = 1'b1; // Expected: {'sum': 134, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b00001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2829,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 134, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100100; b = 8'b10011010; cin = 1'b0; // Expected: {'sum': 62, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100100; b = 8'b10011010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2830,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 62, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b01001111; cin = 1'b1; // Expected: {'sum': 217, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b01001111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2831,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 217, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101111; b = 8'b00011000; cin = 1'b1; // Expected: {'sum': 8, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101111; b = 8'b00011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2832,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 8, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110000; b = 8'b01100110; cin = 1'b0; // Expected: {'sum': 150, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110000; b = 8'b01100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2833,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 150, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111010; b = 8'b10101010; cin = 1'b0; // Expected: {'sum': 164, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111010; b = 8'b10101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2834,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 164, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110110; b = 8'b01000111; cin = 1'b0; // Expected: {'sum': 189, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110110; b = 8'b01000111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2835,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 189, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b10010110; cin = 1'b1; // Expected: {'sum': 36, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b10010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2836,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 36, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101110; b = 8'b00110111; cin = 1'b0; // Expected: {'sum': 101, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101110; b = 8'b00110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2837,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 101, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101111; b = 8'b01010110; cin = 1'b0; // Expected: {'sum': 197, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101111; b = 8'b01010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2838,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 197, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001100; b = 8'b10011100; cin = 1'b1; // Expected: {'sum': 41, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001100; b = 8'b10011100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2839,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 41, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b10000111; cin = 1'b1; // Expected: {'sum': 96, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b10000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2840,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 96, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b00001011; cin = 1'b1; // Expected: {'sum': 127, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b00001011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2841,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 127, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b10011001; cin = 1'b1; // Expected: {'sum': 139, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b10011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2842,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 139, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b11010100; cin = 1'b1; // Expected: {'sum': 218, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b11010100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2843,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 218, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b01110001; cin = 1'b0; // Expected: {'sum': 211, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b01110001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2844,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 211, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b11110101; cin = 1'b1; // Expected: {'sum': 0, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b11110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2845,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b01111000; cin = 1'b1; // Expected: {'sum': 30, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b01111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2846,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 30, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b00000100; cin = 1'b1; // Expected: {'sum': 252, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b00000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2847,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 252, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000101; b = 8'b11110011; cin = 1'b0; // Expected: {'sum': 120, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000101; b = 8'b11110011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2848,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 120, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b11100011; cin = 1'b0; // Expected: {'sum': 232, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b11100011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2849,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 232, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b11011001; cin = 1'b0; // Expected: {'sum': 241, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b11011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2850,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 241, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101000; b = 8'b00011101; cin = 1'b1; // Expected: {'sum': 70, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101000; b = 8'b00011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2851,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 70, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011001; b = 8'b01000001; cin = 1'b1; // Expected: {'sum': 155, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011001; b = 8'b01000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2852,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 155, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b10111010; cin = 1'b1; // Expected: {'sum': 5, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b10111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2853,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 5, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001110; b = 8'b01101111; cin = 1'b1; // Expected: {'sum': 126, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001110; b = 8'b01101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2854,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 126, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b11000010; cin = 1'b1; // Expected: {'sum': 66, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b11000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2855,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 66, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000100; b = 8'b01000111; cin = 1'b1; // Expected: {'sum': 76, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000100; b = 8'b01000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2856,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 76, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110101; b = 8'b00101111; cin = 1'b0; // Expected: {'sum': 228, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110101; b = 8'b00101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2857,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 228, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010101; b = 8'b10010001; cin = 1'b1; // Expected: {'sum': 167, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010101; b = 8'b10010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2858,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 167, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011001; b = 8'b11010000; cin = 1'b0; // Expected: {'sum': 105, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011001; b = 8'b11010000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2859,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 105, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011101; b = 8'b11110110; cin = 1'b1; // Expected: {'sum': 148, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011101; b = 8'b11110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2860,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 148, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b01011110; cin = 1'b0; // Expected: {'sum': 163, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b01011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2861,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 163, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b01101001; cin = 1'b1; // Expected: {'sum': 25, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b01101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2862,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 25, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101010; b = 8'b10101111; cin = 1'b1; // Expected: {'sum': 154, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101010; b = 8'b10101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2863,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 154, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111111; b = 8'b10001010; cin = 1'b0; // Expected: {'sum': 73, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111111; b = 8'b10001010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2864,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 73, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b00111111; cin = 1'b0; // Expected: {'sum': 238, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b00111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2865,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 238, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b11000100; cin = 1'b1; // Expected: {'sum': 70, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b11000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2866,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 70, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b10100110; cin = 1'b0; // Expected: {'sum': 234, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b10100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2867,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 234, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b01100111; cin = 1'b1; // Expected: {'sum': 38, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b01100111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2868,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 38, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100000; b = 8'b01000100; cin = 1'b0; // Expected: {'sum': 36, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100000; b = 8'b01000100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2869,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 36, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010101; b = 8'b11000010; cin = 1'b0; // Expected: {'sum': 215, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010101; b = 8'b11000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2870,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 215, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010000; b = 8'b10111100; cin = 1'b0; // Expected: {'sum': 204, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010000; b = 8'b10111100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2871,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 204, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b01010010; cin = 1'b1; // Expected: {'sum': 169, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b01010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2872,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 169, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b00101000; cin = 1'b0; // Expected: {'sum': 7, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b00101000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2873,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b10010100; cin = 1'b1; // Expected: {'sum': 175, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b10010100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2874,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 175, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b10000101; cin = 1'b0; // Expected: {'sum': 155, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b10000101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2875,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 155, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b01000000; cin = 1'b0; // Expected: {'sum': 188, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b01000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2876,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 188, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001111; b = 8'b10011000; cin = 1'b0; // Expected: {'sum': 231, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001111; b = 8'b10011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2877,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 231, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011101; b = 8'b10010111; cin = 1'b0; // Expected: {'sum': 52, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011101; b = 8'b10010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2878,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 52, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b10001111; cin = 1'b0; // Expected: {'sum': 70, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b10001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2879,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 70, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b00111000; cin = 1'b1; // Expected: {'sum': 55, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b00111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2880,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 55, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b10101001; cin = 1'b1; // Expected: {'sum': 18, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b10101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2881,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 18, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b01100011; cin = 1'b0; // Expected: {'sum': 196, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b01100011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2882,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 196, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b10100100; cin = 1'b0; // Expected: {'sum': 42, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b10100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2883,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 42, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b01110111; cin = 1'b0; // Expected: {'sum': 234, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b01110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2884,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 234, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101100; b = 8'b11100000; cin = 1'b1; // Expected: {'sum': 205, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101100; b = 8'b11100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2885,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 205, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b01010101; cin = 1'b1; // Expected: {'sum': 76, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b01010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2886,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 76, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b00010000; cin = 1'b1; // Expected: {'sum': 75, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b00010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2887,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 75, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100111; b = 8'b10110110; cin = 1'b1; // Expected: {'sum': 222, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100111; b = 8'b10110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2888,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 222, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111111; b = 8'b10101111; cin = 1'b1; // Expected: {'sum': 111, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111111; b = 8'b10101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2889,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 111, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b01110000; cin = 1'b0; // Expected: {'sum': 206, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b01110000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2890,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 206, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b11010111; cin = 1'b0; // Expected: {'sum': 96, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b11010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2891,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 96, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b10100101; cin = 1'b1; // Expected: {'sum': 34, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b10100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2892,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 34, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b01100100; cin = 1'b0; // Expected: {'sum': 191, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b01100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2893,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 191, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b01010010; cin = 1'b1; // Expected: {'sum': 12, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b01010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2894,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000100; b = 8'b00010111; cin = 1'b1; // Expected: {'sum': 28, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000100; b = 8'b00010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2895,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 28, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b10001011; cin = 1'b0; // Expected: {'sum': 254, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b10001011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2896,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 254, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b10100000; cin = 1'b0; // Expected: {'sum': 120, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b10100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2897,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 120, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111011; b = 8'b11011011; cin = 1'b0; // Expected: {'sum': 150, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111011; b = 8'b11011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2898,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 150, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b10101110; cin = 1'b0; // Expected: {'sum': 242, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b10101110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2899,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 242, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b01101000; cin = 1'b1; // Expected: {'sum': 242, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b01101000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2900,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 242, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111010; b = 8'b00111010; cin = 1'b1; // Expected: {'sum': 53, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111010; b = 8'b00111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2901,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 53, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110111; b = 8'b11011101; cin = 1'b1; // Expected: {'sum': 21, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110111; b = 8'b11011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2902,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 21, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b00001010; cin = 1'b1; // Expected: {'sum': 30, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b00001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2903,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 30, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b01100001; cin = 1'b1; // Expected: {'sum': 192, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b01100001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2904,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 192, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b01100000; cin = 1'b0; // Expected: {'sum': 63, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b01100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2905,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 63, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110111; b = 8'b01010110; cin = 1'b0; // Expected: {'sum': 141, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110111; b = 8'b01010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2906,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 141, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b00000000; cin = 1'b0; // Expected: {'sum': 41, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b00000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2907,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 41, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b01100001; cin = 1'b0; // Expected: {'sum': 49, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b01100001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2908,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 49, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b00111011; cin = 1'b0; // Expected: {'sum': 247, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b00111011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2909,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 247, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000011; b = 8'b00001011; cin = 1'b0; // Expected: {'sum': 206, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000011; b = 8'b00001011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2910,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 206, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010010; b = 8'b10110010; cin = 1'b0; // Expected: {'sum': 4, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010010; b = 8'b10110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2911,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b11101000; cin = 1'b0; // Expected: {'sum': 118, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b11101000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2912,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 118, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b01011011; cin = 1'b0; // Expected: {'sum': 41, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b01011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2913,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 41, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011010; b = 8'b10001100; cin = 1'b1; // Expected: {'sum': 103, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011010; b = 8'b10001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2914,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 103, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b10011110; cin = 1'b0; // Expected: {'sum': 36, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b10011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2915,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 36, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b11000100; cin = 1'b1; // Expected: {'sum': 71, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b11000100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2916,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 71, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b01000110; cin = 1'b1; // Expected: {'sum': 178, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b01000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2917,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 178, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b10100000; cin = 1'b1; // Expected: {'sum': 230, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b10100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2918,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 230, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001100; b = 8'b10010100; cin = 1'b0; // Expected: {'sum': 160, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001100; b = 8'b10010100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2919,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 160, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b01011000; cin = 1'b1; // Expected: {'sum': 156, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b01011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2920,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 156, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100100; b = 8'b11011111; cin = 1'b1; // Expected: {'sum': 132, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100100; b = 8'b11011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2921,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 132, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111000; b = 8'b01010001; cin = 1'b0; // Expected: {'sum': 137, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111000; b = 8'b01010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2922,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 137, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001101; b = 8'b00011101; cin = 1'b1; // Expected: {'sum': 235, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001101; b = 8'b00011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2923,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 235, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b01000000; cin = 1'b0; // Expected: {'sum': 124, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b01000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2924,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 124, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101000; b = 8'b01111100; cin = 1'b0; // Expected: {'sum': 164, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101000; b = 8'b01111100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2925,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 164, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b01111010; cin = 1'b0; // Expected: {'sum': 29, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b01111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2926,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 29, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010000; b = 8'b10100011; cin = 1'b0; // Expected: {'sum': 179, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010000; b = 8'b10100011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2927,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 179, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b10001001; cin = 1'b1; // Expected: {'sum': 133, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b10001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2928,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 133, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100111; b = 8'b00011100; cin = 1'b0; // Expected: {'sum': 131, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100111; b = 8'b00011100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2929,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 131, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111001; b = 8'b00001001; cin = 1'b1; // Expected: {'sum': 67, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111001; b = 8'b00001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2930,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 67, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b00000100; cin = 1'b0; // Expected: {'sum': 192, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b00000100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2931,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 192, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b01110001; cin = 1'b1; // Expected: {'sum': 220, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b01110001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2932,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 220, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b10001100; cin = 1'b0; // Expected: {'sum': 171, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b10001100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2933,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 171, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b01001100; cin = 1'b0; // Expected: {'sum': 107, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b01001100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2934,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 107, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b10101110; cin = 1'b0; // Expected: {'sum': 162, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b10101110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2935,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 162, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001011; b = 8'b00101100; cin = 1'b0; // Expected: {'sum': 55, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001011; b = 8'b00101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2936,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 55, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b10010001; cin = 1'b1; // Expected: {'sum': 134, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b10010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2937,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 134, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011110; b = 8'b01111110; cin = 1'b0; // Expected: {'sum': 92, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011110; b = 8'b01111110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2938,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 92, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b01111010; cin = 1'b1; // Expected: {'sum': 254, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b01111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2939,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 254, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000111; b = 8'b00111111; cin = 1'b0; // Expected: {'sum': 198, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000111; b = 8'b00111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2940,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 198, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101110; b = 8'b00110101; cin = 1'b1; // Expected: {'sum': 228, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101110; b = 8'b00110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2941,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 228, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101100; b = 8'b01101100; cin = 1'b1; // Expected: {'sum': 25, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101100; b = 8'b01101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2942,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 25, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b10110011; cin = 1'b0; // Expected: {'sum': 210, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b10110011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2943,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 210, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b11101011; cin = 1'b0; // Expected: {'sum': 73, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b11101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2944,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 73, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b10110010; cin = 1'b0; // Expected: {'sum': 46, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b10110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2945,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 46, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010001; b = 8'b01111101; cin = 1'b1; // Expected: {'sum': 79, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010001; b = 8'b01111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2946,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 79, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b11000011; cin = 1'b1; // Expected: {'sum': 86, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b11000011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2947,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 86, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b10010100; cin = 1'b0; // Expected: {'sum': 22, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b10010100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2948,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 22, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b01110110; cin = 1'b1; // Expected: {'sum': 71, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b01110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2949,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 71, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b00100111; cin = 1'b1; // Expected: {'sum': 201, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b00100111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2950,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 201, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b11110101; cin = 1'b0; // Expected: {'sum': 191, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b11110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2951,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 191, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b10000011; cin = 1'b0; // Expected: {'sum': 212, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b10000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2952,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 212, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001111; b = 8'b00000000; cin = 1'b1; // Expected: {'sum': 80, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001111; b = 8'b00000000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2953,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 80, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101100; b = 8'b01111110; cin = 1'b0; // Expected: {'sum': 106, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101100; b = 8'b01111110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2954,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 106, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b11011010; cin = 1'b1; // Expected: {'sum': 64, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b11011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2955,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 64, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110011; b = 8'b00000000; cin = 1'b1; // Expected: {'sum': 180, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110011; b = 8'b00000000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2956,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 180, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b10011111; cin = 1'b1; // Expected: {'sum': 228, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b10011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2957,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 228, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b00100001; cin = 1'b1; // Expected: {'sum': 194, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b00100001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2958,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 194, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100000; b = 8'b01000111; cin = 1'b0; // Expected: {'sum': 167, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100000; b = 8'b01000111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2959,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 167, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b00101011; cin = 1'b1; // Expected: {'sum': 34, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b00101011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2960,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 34, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111011; b = 8'b00100011; cin = 1'b0; // Expected: {'sum': 158, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111011; b = 8'b00100011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2961,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 158, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b11011110; cin = 1'b0; // Expected: {'sum': 97, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b11011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2962,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 97, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b01011101; cin = 1'b1; // Expected: {'sum': 92, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b01011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2963,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 92, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100010; b = 8'b01111001; cin = 1'b1; // Expected: {'sum': 92, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100010; b = 8'b01111001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2964,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 92, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b01110001; cin = 1'b1; // Expected: {'sum': 8, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b01110001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2965,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 8, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b10111011; cin = 1'b1; // Expected: {'sum': 81, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b10111011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2966,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 81, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110110; b = 8'b01000011; cin = 1'b1; // Expected: {'sum': 186, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110110; b = 8'b01000011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2967,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 186, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b01011110; cin = 1'b0; // Expected: {'sum': 54, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b01011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2968,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 54, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b01000101; cin = 1'b1; // Expected: {'sum': 16, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b01000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2969,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 16, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b11100000; cin = 1'b0; // Expected: {'sum': 157, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b11100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2970,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 157, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b10101000; cin = 1'b1; // Expected: {'sum': 55, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b10101000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2971,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 55, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001101; b = 8'b10000010; cin = 1'b1; // Expected: {'sum': 144, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001101; b = 8'b10000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2972,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 144, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100100; b = 8'b10011001; cin = 1'b0; // Expected: {'sum': 61, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100100; b = 8'b10011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2973,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 61, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b11110001; cin = 1'b1; // Expected: {'sum': 176, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b11110001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2974,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 176, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000000; b = 8'b01111001; cin = 1'b1; // Expected: {'sum': 250, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000000; b = 8'b01111001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2975,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 250, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b11101011; cin = 1'b0; // Expected: {'sum': 148, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b11101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2976,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 148, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100011; b = 8'b01001100; cin = 1'b0; // Expected: {'sum': 47, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100011; b = 8'b01001100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2977,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 47, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b11010101; cin = 1'b1; // Expected: {'sum': 183, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b11010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2978,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 183, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b11111100; cin = 1'b0; // Expected: {'sum': 184, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b11111100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2979,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 184, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b00100000; cin = 1'b1; // Expected: {'sum': 119, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b00100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2980,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 119, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b10010101; cin = 1'b0; // Expected: {'sum': 106, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b10010101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2981,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 106, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001001; b = 8'b11111110; cin = 1'b1; // Expected: {'sum': 72, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001001; b = 8'b11111110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2982,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 72, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b01001110; cin = 1'b0; // Expected: {'sum': 171, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b01001110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2983,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 171, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b11000111; cin = 1'b1; // Expected: {'sum': 35, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b11000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2984,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 35, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b10101111; cin = 1'b0; // Expected: {'sum': 198, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b10101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2985,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 198, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010011; b = 8'b01100100; cin = 1'b0; // Expected: {'sum': 247, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010011; b = 8'b01100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2986,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 247, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010101; b = 8'b00011000; cin = 1'b1; // Expected: {'sum': 46, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010101; b = 8'b00011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2987,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 46, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b11101110; cin = 1'b0; // Expected: {'sum': 157, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b11101110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2988,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 157, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b11001000; cin = 1'b1; // Expected: {'sum': 245, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b11001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2989,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 245, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b00101101; cin = 1'b1; // Expected: {'sum': 140, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b00101101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2990,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 140, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010010; b = 8'b01100111; cin = 1'b0; // Expected: {'sum': 185, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010010; b = 8'b01100111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2991,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 185, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111011; b = 8'b11001101; cin = 1'b0; // Expected: {'sum': 8, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111011; b = 8'b11001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2992,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 8, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b01001111; cin = 1'b0; // Expected: {'sum': 12, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b01001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2993,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b01010110; cin = 1'b0; // Expected: {'sum': 120, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b01010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2994,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 120, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b01100111; cin = 1'b0; // Expected: {'sum': 234, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b01100111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2995,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 234, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b01110101; cin = 1'b0; // Expected: {'sum': 232, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b01110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2996,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 232, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b10010110; cin = 1'b1; // Expected: {'sum': 203, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b10010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2997,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 203, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b10010000; cin = 1'b0; // Expected: {'sum': 188, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b10010000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2998,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 188, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b01100111; cin = 1'b0; // Expected: {'sum': 133, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b01100111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2999,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 133, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b00010100; cin = 1'b1; // Expected: {'sum': 127, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b00010100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3000,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 127, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b00100000; cin = 1'b1; // Expected: {'sum': 160, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b00100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3001,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 160, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011100; b = 8'b11101100; cin = 1'b1; // Expected: {'sum': 201, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011100; b = 8'b11101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3002,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 201, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b10110110; cin = 1'b1; // Expected: {'sum': 31, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b10110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3003,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 31, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b01100100; cin = 1'b0; // Expected: {'sum': 231, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b01100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3004,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 231, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b01101110; cin = 1'b1; // Expected: {'sum': 180, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b01101110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3005,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 180, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b10000111; cin = 1'b1; // Expected: {'sum': 171, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b10000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3006,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 171, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b00011110; cin = 1'b1; // Expected: {'sum': 155, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b00011110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3007,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 155, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b01000001; cin = 1'b0; // Expected: {'sum': 251, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b01000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3008,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 251, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b00011101; cin = 1'b0; // Expected: {'sum': 73, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b00011101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3009,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 73, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b11011010; cin = 1'b1; // Expected: {'sum': 30, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b11011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3010,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 30, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001111; b = 8'b00110101; cin = 1'b1; // Expected: {'sum': 133, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001111; b = 8'b00110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3011,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 133, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b11001110; cin = 1'b1; // Expected: {'sum': 158, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b11001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3012,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 158, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b00011000; cin = 1'b0; // Expected: {'sum': 92, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b00011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3013,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 92, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010001; b = 8'b00111011; cin = 1'b1; // Expected: {'sum': 13, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010001; b = 8'b00111011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3014,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 13, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001001; b = 8'b01000010; cin = 1'b1; // Expected: {'sum': 12, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001001; b = 8'b01000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3015,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b11000011; cin = 1'b0; // Expected: {'sum': 37, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b11000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3016,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 37, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b01111010; cin = 1'b0; // Expected: {'sum': 18, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b01111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3017,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 18, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b11111000; cin = 1'b1; // Expected: {'sum': 228, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b11111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3018,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 228, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b01001100; cin = 1'b1; // Expected: {'sum': 10, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b01001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3019,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001000; b = 8'b11110111; cin = 1'b1; // Expected: {'sum': 64, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001000; b = 8'b11110111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3020,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 64, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b10110110; cin = 1'b0; // Expected: {'sum': 142, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b10110110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3021,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 142, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b10011111; cin = 1'b1; // Expected: {'sum': 197, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b10011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3022,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 197, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101100; b = 8'b00100001; cin = 1'b1; // Expected: {'sum': 14, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101100; b = 8'b00100001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3023,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b00010000; cin = 1'b1; // Expected: {'sum': 211, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b00010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3024,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 211, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b01000010; cin = 1'b0; // Expected: {'sum': 157, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b01000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3025,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 157, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b01111010; cin = 1'b0; // Expected: {'sum': 7, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b01111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3026,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010101; b = 8'b11011101; cin = 1'b0; // Expected: {'sum': 50, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010101; b = 8'b11011101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3027,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 50, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b00101110; cin = 1'b0; // Expected: {'sum': 7, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b00101110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3028,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b11000001; cin = 1'b0; // Expected: {'sum': 129, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b11000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3029,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 129, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011111; b = 8'b10110010; cin = 1'b0; // Expected: {'sum': 81, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011111; b = 8'b10110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3030,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 81, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b10101100; cin = 1'b1; // Expected: {'sum': 227, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b10101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3031,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 227, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b10000101; cin = 1'b1; // Expected: {'sum': 141, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b10000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3032,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 141, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000111; b = 8'b00101000; cin = 1'b1; // Expected: {'sum': 176, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000111; b = 8'b00101000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3033,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 176, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100100; b = 8'b11010101; cin = 1'b1; // Expected: {'sum': 122, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100100; b = 8'b11010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3034,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 122, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b00110100; cin = 1'b1; // Expected: {'sum': 242, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b00110100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3035,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 242, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b01110100; cin = 1'b0; // Expected: {'sum': 123, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b01110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3036,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 123, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b00010110; cin = 1'b0; // Expected: {'sum': 251, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b00010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3037,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 251, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b01001100; cin = 1'b1; // Expected: {'sum': 255, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b01001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3038,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 255, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b11110001; cin = 1'b0; // Expected: {'sum': 228, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b11110001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3039,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 228, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111000; b = 8'b10011000; cin = 1'b0; // Expected: {'sum': 208, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111000; b = 8'b10011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3040,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 208, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001101; b = 8'b11000101; cin = 1'b0; // Expected: {'sum': 210, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001101; b = 8'b11000101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3041,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 210, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b00100010; cin = 1'b1; // Expected: {'sum': 166, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b00100010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3042,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 166, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b01100011; cin = 1'b0; // Expected: {'sum': 208, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b01100011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3043,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 208, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b01010110; cin = 1'b1; // Expected: {'sum': 214, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b01010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3044,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 214, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011101; b = 8'b01011100; cin = 1'b1; // Expected: {'sum': 250, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011101; b = 8'b01011100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3045,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 250, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111000; b = 8'b11000000; cin = 1'b0; // Expected: {'sum': 248, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111000; b = 8'b11000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3046,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 248, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001100; b = 8'b11110101; cin = 1'b1; // Expected: {'sum': 194, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001100; b = 8'b11110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3047,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 194, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b10001111; cin = 1'b0; // Expected: {'sum': 148, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b10001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3048,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 148, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b01101010; cin = 1'b1; // Expected: {'sum': 176, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b01101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3049,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 176, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011111; b = 8'b01000011; cin = 1'b0; // Expected: {'sum': 162, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011111; b = 8'b01000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3050,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 162, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001011; b = 8'b10001011; cin = 1'b1; // Expected: {'sum': 215, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001011; b = 8'b10001011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3051,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 215, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b00111101; cin = 1'b1; // Expected: {'sum': 31, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b00111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3052,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 31, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b00101001; cin = 1'b0; // Expected: {'sum': 117, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b00101001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3053,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 117, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b01111010; cin = 1'b0; // Expected: {'sum': 34, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b01111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3054,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 34, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b10111011; cin = 1'b1; // Expected: {'sum': 59, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b10111011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3055,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 59, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b11000000; cin = 1'b1; // Expected: {'sum': 217, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b11000000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3056,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 217, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b01111100; cin = 1'b1; // Expected: {'sum': 63, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b01111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3057,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 63, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110101; b = 8'b01010100; cin = 1'b1; // Expected: {'sum': 138, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110101; b = 8'b01010100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3058,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 138, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001011; b = 8'b11000101; cin = 1'b0; // Expected: {'sum': 208, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001011; b = 8'b11000101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3059,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 208, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b10110101; cin = 1'b0; // Expected: {'sum': 255, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b10110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3060,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 255, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100111; b = 8'b10101110; cin = 1'b1; // Expected: {'sum': 86, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100111; b = 8'b10101110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3061,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 86, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b00110010; cin = 1'b1; // Expected: {'sum': 209, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b00110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3062,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 209, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100001; b = 8'b11010101; cin = 1'b0; // Expected: {'sum': 246, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100001; b = 8'b11010101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3063,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 246, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010100; b = 8'b00100101; cin = 1'b0; // Expected: {'sum': 249, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010100; b = 8'b00100101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3064,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 249, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b01010111; cin = 1'b1; // Expected: {'sum': 90, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b01010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3065,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 90, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011111; b = 8'b11110010; cin = 1'b1; // Expected: {'sum': 146, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011111; b = 8'b11110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3066,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 146, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b01100010; cin = 1'b1; // Expected: {'sum': 50, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b01100010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3067,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 50, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b01011100; cin = 1'b0; // Expected: {'sum': 52, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b01011100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3068,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 52, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b00111111; cin = 1'b1; // Expected: {'sum': 114, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b00111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3069,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 114, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b01110000; cin = 1'b1; // Expected: {'sum': 235, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b01110000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3070,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 235, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b10010010; cin = 1'b1; // Expected: {'sum': 147, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b10010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3071,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 147, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011010; b = 8'b01110100; cin = 1'b0; // Expected: {'sum': 14, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011010; b = 8'b01110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3072,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001010; b = 8'b10100110; cin = 1'b0; // Expected: {'sum': 48, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001010; b = 8'b10100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3073,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 48, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b11011100; cin = 1'b0; // Expected: {'sum': 142, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b11011100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3074,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 142, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b01101001; cin = 1'b1; // Expected: {'sum': 243, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b01101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3075,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 243, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b11110111; cin = 1'b0; // Expected: {'sum': 132, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b11110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3076,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 132, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b01011000; cin = 1'b1; // Expected: {'sum': 48, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b01011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3077,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 48, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b11110010; cin = 1'b0; // Expected: {'sum': 240, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b11110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3078,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 240, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101000; b = 8'b01010111; cin = 1'b0; // Expected: {'sum': 127, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101000; b = 8'b01010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3079,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 127, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001111; b = 8'b10100011; cin = 1'b0; // Expected: {'sum': 242, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001111; b = 8'b10100011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3080,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 242, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001001; b = 8'b10000111; cin = 1'b0; // Expected: {'sum': 80, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001001; b = 8'b10000111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3081,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 80, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b01110011; cin = 1'b0; // Expected: {'sum': 189, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b01110011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3082,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 189, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100110; b = 8'b01010001; cin = 1'b0; // Expected: {'sum': 55, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100110; b = 8'b01010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3083,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 55, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b11000110; cin = 1'b1; // Expected: {'sum': 253, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b11000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3084,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 253, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b00101100; cin = 1'b0; // Expected: {'sum': 240, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b00101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3085,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 240, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b00000101; cin = 1'b0; // Expected: {'sum': 59, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b00000101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3086,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 59, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110100; b = 8'b00010101; cin = 1'b0; // Expected: {'sum': 137, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110100; b = 8'b00010101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3087,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 137, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101010; b = 8'b01101010; cin = 1'b0; // Expected: {'sum': 20, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101010; b = 8'b01101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3088,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 20, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100000; b = 8'b10011110; cin = 1'b0; // Expected: {'sum': 254, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100000; b = 8'b10011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3089,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 254, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b01100101; cin = 1'b0; // Expected: {'sum': 124, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b01100101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3090,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 124, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b11110111; cin = 1'b0; // Expected: {'sum': 112, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b11110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3091,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 112, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010100; b = 8'b00011101; cin = 1'b1; // Expected: {'sum': 114, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010100; b = 8'b00011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3092,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 114, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b01011100; cin = 1'b0; // Expected: {'sum': 46, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b01011100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3093,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 46, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b00111100; cin = 1'b0; // Expected: {'sum': 69, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b00111100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3094,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 69, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000110; b = 8'b10011011; cin = 1'b1; // Expected: {'sum': 162, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000110; b = 8'b10011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3095,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 162, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111011; b = 8'b01111000; cin = 1'b1; // Expected: {'sum': 52, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111011; b = 8'b01111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3096,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 52, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b11111010; cin = 1'b1; // Expected: {'sum': 208, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b11111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3097,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 208, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b10011111; cin = 1'b1; // Expected: {'sum': 226, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b10011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3098,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 226, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000111; b = 8'b01110000; cin = 1'b0; // Expected: {'sum': 55, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000111; b = 8'b01110000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3099,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 55, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b00001010; cin = 1'b0; // Expected: {'sum': 32, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b00001010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3100,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 32, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b10010101; cin = 1'b1; // Expected: {'sum': 117, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b10010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3101,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 117, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b00000000; cin = 1'b0; // Expected: {'sum': 132, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b00000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3102,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 132, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b00000101; cin = 1'b1; // Expected: {'sum': 41, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b00000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3103,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 41, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111001; b = 8'b01001011; cin = 1'b1; // Expected: {'sum': 133, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111001; b = 8'b01001011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3104,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 133, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b10011101; cin = 1'b1; // Expected: {'sum': 34, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b10011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3105,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 34, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010010; b = 8'b11001001; cin = 1'b0; // Expected: {'sum': 219, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010010; b = 8'b11001001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3106,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 219, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001111; b = 8'b10010100; cin = 1'b0; // Expected: {'sum': 163, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001111; b = 8'b10010100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3107,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 163, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b11011101; cin = 1'b1; // Expected: {'sum': 7, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b11011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3108,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b01001100; cin = 1'b1; // Expected: {'sum': 246, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b01001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3109,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 246, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b00010111; cin = 1'b0; // Expected: {'sum': 147, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b00010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3110,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 147, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b10110101; cin = 1'b1; // Expected: {'sum': 248, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b10110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3111,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 248, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b00001101; cin = 1'b1; // Expected: {'sum': 200, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b00001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3112,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 200, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b01100110; cin = 1'b1; // Expected: {'sum': 16, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b01100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3113,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 16, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b11000101; cin = 1'b1; // Expected: {'sum': 11, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b11000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3114,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 11, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b01001101; cin = 1'b1; // Expected: {'sum': 164, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b01001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3115,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 164, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101111; b = 8'b01101000; cin = 1'b1; // Expected: {'sum': 88, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101111; b = 8'b01101000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3116,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 88, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b01001001; cin = 1'b0; // Expected: {'sum': 170, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b01001001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3117,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 170, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001011; b = 8'b10001000; cin = 1'b0; // Expected: {'sum': 211, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001011; b = 8'b10001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3118,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 211, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001100; b = 8'b10001101; cin = 1'b1; // Expected: {'sum': 90, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001100; b = 8'b10001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3119,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 90, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101111; b = 8'b01001001; cin = 1'b0; // Expected: {'sum': 120, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101111; b = 8'b01001001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3120,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 120, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000111; b = 8'b00100100; cin = 1'b1; // Expected: {'sum': 172, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000111; b = 8'b00100100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3121,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 172, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110000; b = 8'b10101101; cin = 1'b1; // Expected: {'sum': 30, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110000; b = 8'b10101101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3122,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 30, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011101; b = 8'b10001000; cin = 1'b0; // Expected: {'sum': 101, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011101; b = 8'b10001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3123,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 101, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101010; b = 8'b01010010; cin = 1'b0; // Expected: {'sum': 124, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101010; b = 8'b01010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3124,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 124, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b11100111; cin = 1'b0; // Expected: {'sum': 82, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b11100111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3125,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 82, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011101; b = 8'b10000001; cin = 1'b0; // Expected: {'sum': 94, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011101; b = 8'b10000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3126,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 94, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b01010110; cin = 1'b0; // Expected: {'sum': 186, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b01010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3127,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 186, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b10010110; cin = 1'b0; // Expected: {'sum': 96, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b10010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3128,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 96, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b01001001; cin = 1'b1; // Expected: {'sum': 69, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b01001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3129,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 69, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b01010110; cin = 1'b1; // Expected: {'sum': 138, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b01010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3130,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 138, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010011; b = 8'b11100000; cin = 1'b0; // Expected: {'sum': 179, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010011; b = 8'b11100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3131,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 179, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101001; b = 8'b11000110; cin = 1'b1; // Expected: {'sum': 48, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101001; b = 8'b11000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3132,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 48, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100100; b = 8'b01001010; cin = 1'b0; // Expected: {'sum': 238, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100100; b = 8'b01001010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3133,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 238, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b00000111; cin = 1'b0; // Expected: {'sum': 159, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b00000111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3134,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 159, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010010; b = 8'b11011010; cin = 1'b1; // Expected: {'sum': 237, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010010; b = 8'b11011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3135,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 237, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b01011000; cin = 1'b1; // Expected: {'sum': 157, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b01011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3136,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 157, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010111; b = 8'b10010101; cin = 1'b0; // Expected: {'sum': 236, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010111; b = 8'b10010101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3137,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 236, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101011; b = 8'b10011001; cin = 1'b0; // Expected: {'sum': 196, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101011; b = 8'b10011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3138,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 196, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b01010011; cin = 1'b0; // Expected: {'sum': 10, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b01010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3139,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b00001110; cin = 1'b0; // Expected: {'sum': 49, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b00001110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3140,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 49, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b00101010; cin = 1'b0; // Expected: {'sum': 72, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b00101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3141,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 72, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b10100001; cin = 1'b1; // Expected: {'sum': 36, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b10100001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3142,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 36, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b00100011; cin = 1'b0; // Expected: {'sum': 111, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b00100011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3143,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 111, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010011; b = 8'b01011101; cin = 1'b1; // Expected: {'sum': 241, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010011; b = 8'b01011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3144,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 241, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b00110111; cin = 1'b1; // Expected: {'sum': 202, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b00110111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3145,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 202, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011010; b = 8'b11110110; cin = 1'b0; // Expected: {'sum': 80, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011010; b = 8'b11110110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3146,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 80, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b11001010; cin = 1'b1; // Expected: {'sum': 99, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b11001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3147,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 99, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b01010100; cin = 1'b0; // Expected: {'sum': 20, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b01010100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3148,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 20, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b11000001; cin = 1'b0; // Expected: {'sum': 183, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b11000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3149,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 183, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b10001010; cin = 1'b0; // Expected: {'sum': 236, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b10001010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3150,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 236, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100111; b = 8'b00111110; cin = 1'b1; // Expected: {'sum': 38, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100111; b = 8'b00111110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3151,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 38, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b00010000; cin = 1'b0; // Expected: {'sum': 185, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b00010000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3152,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 185, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100111; b = 8'b01111000; cin = 1'b1; // Expected: {'sum': 160, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100111; b = 8'b01111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3153,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 160, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b01010001; cin = 1'b0; // Expected: {'sum': 103, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b01010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3154,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 103, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b00001110; cin = 1'b1; // Expected: {'sum': 124, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b00001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3155,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 124, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b01100100; cin = 1'b1; // Expected: {'sum': 168, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b01100100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3156,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 168, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b11110000; cin = 1'b0; // Expected: {'sum': 227, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b11110000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3157,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 227, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001101; b = 8'b11001001; cin = 1'b0; // Expected: {'sum': 150, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001101; b = 8'b11001001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3158,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 150, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000110; b = 8'b10010000; cin = 1'b1; // Expected: {'sum': 87, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000110; b = 8'b10010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3159,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 87, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b11111010; cin = 1'b0; // Expected: {'sum': 4, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b11111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3160,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101110; b = 8'b00110010; cin = 1'b1; // Expected: {'sum': 97, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101110; b = 8'b00110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3161,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 97, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b00001101; cin = 1'b1; // Expected: {'sum': 136, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b00001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3162,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 136, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b11111110; cin = 1'b0; // Expected: {'sum': 17, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b11111110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3163,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 17, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110101; b = 8'b00111100; cin = 1'b1; // Expected: {'sum': 114, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110101; b = 8'b00111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3164,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 114, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b10010111; cin = 1'b1; // Expected: {'sum': 54, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b10010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3165,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 54, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100110; b = 8'b01001110; cin = 1'b1; // Expected: {'sum': 53, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100110; b = 8'b01001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3166,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 53, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b00111010; cin = 1'b1; // Expected: {'sum': 156, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b00111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3167,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 156, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100000; b = 8'b01001110; cin = 1'b0; // Expected: {'sum': 174, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100000; b = 8'b01001110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3168,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 174, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b00001000; cin = 1'b0; // Expected: {'sum': 176, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b00001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3169,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 176, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b00000101; cin = 1'b1; // Expected: {'sum': 244, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b00000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3170,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 244, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110101; b = 8'b11110100; cin = 1'b0; // Expected: {'sum': 169, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110101; b = 8'b11110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3171,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 169, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101001; b = 8'b11001101; cin = 1'b0; // Expected: {'sum': 182, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101001; b = 8'b11001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3172,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 182, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b10111010; cin = 1'b1; // Expected: {'sum': 121, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b10111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3173,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 121, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001111; b = 8'b10011111; cin = 1'b1; // Expected: {'sum': 175, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001111; b = 8'b10011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3174,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 175, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011010; b = 8'b10011010; cin = 1'b1; // Expected: {'sum': 53, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011010; b = 8'b10011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3175,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 53, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011001; b = 8'b00000010; cin = 1'b0; // Expected: {'sum': 91, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011001; b = 8'b00000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3176,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 91, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011001; b = 8'b01100000; cin = 1'b1; // Expected: {'sum': 122, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011001; b = 8'b01100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3177,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 122, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111001; b = 8'b11111010; cin = 1'b0; // Expected: {'sum': 51, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111001; b = 8'b11111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3178,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 51, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b10001110; cin = 1'b0; // Expected: {'sum': 240, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b10001110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3179,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 240, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b10001000; cin = 1'b1; // Expected: {'sum': 49, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b10001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3180,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 49, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100011; b = 8'b10001001; cin = 1'b1; // Expected: {'sum': 109, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100011; b = 8'b10001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3181,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 109, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b01001001; cin = 1'b0; // Expected: {'sum': 215, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b01001001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3182,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 215, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b10011111; cin = 1'b1; // Expected: {'sum': 86, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b10011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3183,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 86, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b11001010; cin = 1'b1; // Expected: {'sum': 97, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b11001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3184,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 97, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b00010011; cin = 1'b0; // Expected: {'sum': 146, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b00010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3185,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 146, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b11001100; cin = 1'b1; // Expected: {'sum': 213, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b11001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3186,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 213, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101011; b = 8'b01000010; cin = 1'b1; // Expected: {'sum': 110, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101011; b = 8'b01000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3187,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 110, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b10101010; cin = 1'b0; // Expected: {'sum': 99, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b10101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3188,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 99, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011001; b = 8'b11101111; cin = 1'b1; // Expected: {'sum': 73, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011001; b = 8'b11101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3189,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 73, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b00000000; cin = 1'b1; // Expected: {'sum': 207, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b00000000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3190,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 207, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011101; b = 8'b01110000; cin = 1'b1; // Expected: {'sum': 78, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011101; b = 8'b01110000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3191,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 78, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b11001100; cin = 1'b0; // Expected: {'sum': 16, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b11001100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3192,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 16, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101101; b = 8'b10110000; cin = 1'b0; // Expected: {'sum': 93, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101101; b = 8'b10110000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3193,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 93, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b11100011; cin = 1'b0; // Expected: {'sum': 165, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b11100011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3194,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 165, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b10110100; cin = 1'b0; // Expected: {'sum': 116, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b10110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3195,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 116, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b10110011; cin = 1'b0; // Expected: {'sum': 161, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b10110011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3196,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 161, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b00010111; cin = 1'b0; // Expected: {'sum': 92, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b00010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3197,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 92, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b01111010; cin = 1'b1; // Expected: {'sum': 96, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b01111010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3198,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 96, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011010; b = 8'b00011100; cin = 1'b1; // Expected: {'sum': 247, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011010; b = 8'b00011100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3199,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 247, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b11000011; cin = 1'b0; // Expected: {'sum': 133, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b11000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3200,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 133, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010100; b = 8'b11000111; cin = 1'b0; // Expected: {'sum': 219, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010100; b = 8'b11000111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3201,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 219, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b01000101; cin = 1'b0; // Expected: {'sum': 98, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b01000101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3202,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 98, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b01100100; cin = 1'b0; // Expected: {'sum': 13, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b01100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3203,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 13, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b10000011; cin = 1'b0; // Expected: {'sum': 168, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b10000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3204,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 168, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b11001001; cin = 1'b0; // Expected: {'sum': 105, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b11001001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3205,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 105, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b11001100; cin = 1'b0; // Expected: {'sum': 99, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b11001100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3206,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 99, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b00010010; cin = 1'b0; // Expected: {'sum': 118, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b00010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3207,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 118, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b01111010; cin = 1'b0; // Expected: {'sum': 120, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b01111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3208,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 120, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b01010010; cin = 1'b0; // Expected: {'sum': 234, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b01010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3209,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 234, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101001; b = 8'b10110100; cin = 1'b0; // Expected: {'sum': 157, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101001; b = 8'b10110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3210,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 157, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010011; b = 8'b00011101; cin = 1'b1; // Expected: {'sum': 177, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010011; b = 8'b00011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3211,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 177, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101111; b = 8'b10101100; cin = 1'b1; // Expected: {'sum': 28, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101111; b = 8'b10101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3212,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 28, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b11101011; cin = 1'b1; // Expected: {'sum': 231, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b11101011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3213,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 231, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b10111100; cin = 1'b1; // Expected: {'sum': 139, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b10111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3214,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 139, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011010; b = 8'b11010010; cin = 1'b1; // Expected: {'sum': 109, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011010; b = 8'b11010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3215,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 109, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011111; b = 8'b10111100; cin = 1'b1; // Expected: {'sum': 28, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011111; b = 8'b10111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3216,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 28, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b11010010; cin = 1'b1; // Expected: {'sum': 111, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b11010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3217,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 111, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b00100000; cin = 1'b0; // Expected: {'sum': 55, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b00100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3218,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 55, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101001; b = 8'b10111101; cin = 1'b1; // Expected: {'sum': 39, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101001; b = 8'b10111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3219,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 39, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101111; b = 8'b11110110; cin = 1'b0; // Expected: {'sum': 37, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101111; b = 8'b11110110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3220,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 37, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b00100101; cin = 1'b0; // Expected: {'sum': 131, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b00100101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3221,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 131, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b01100000; cin = 1'b1; // Expected: {'sum': 147, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b01100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3222,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 147, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111111; b = 8'b11011101; cin = 1'b0; // Expected: {'sum': 156, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111111; b = 8'b11011101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3223,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 156, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b10011111; cin = 1'b1; // Expected: {'sum': 93, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b10011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3224,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 93, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b00011101; cin = 1'b0; // Expected: {'sum': 20, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b00011101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3225,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 20, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b10001011; cin = 1'b0; // Expected: {'sum': 132, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b10001011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3226,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 132, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b11100010; cin = 1'b0; // Expected: {'sum': 47, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b11100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3227,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 47, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b10111001; cin = 1'b1; // Expected: {'sum': 182, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b10111001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3228,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 182, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100000; b = 8'b01001110; cin = 1'b1; // Expected: {'sum': 47, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100000; b = 8'b01001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3229,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 47, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101010; b = 8'b01111111; cin = 1'b0; // Expected: {'sum': 41, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101010; b = 8'b01111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3230,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 41, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b01000011; cin = 1'b0; // Expected: {'sum': 242, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b01000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3231,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 242, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b00100000; cin = 1'b1; // Expected: {'sum': 87, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b00100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3232,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 87, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b01100111; cin = 1'b1; // Expected: {'sum': 243, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b01100111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3233,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 243, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b10001000; cin = 1'b0; // Expected: {'sum': 181, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b10001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3234,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 181, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010001; b = 8'b10010110; cin = 1'b1; // Expected: {'sum': 104, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010001; b = 8'b10010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3235,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 104, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b11100011; cin = 1'b1; // Expected: {'sum': 63, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b11100011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3236,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 63, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b00101100; cin = 1'b0; // Expected: {'sum': 125, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b00101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3237,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 125, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110001; b = 8'b10010111; cin = 1'b1; // Expected: {'sum': 201, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110001; b = 8'b10010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3238,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 201, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b00000001; cin = 1'b1; // Expected: {'sum': 221, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b00000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3239,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 221, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111011; b = 8'b01000110; cin = 1'b0; // Expected: {'sum': 129, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111011; b = 8'b01000110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3240,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 129, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b10011111; cin = 1'b0; // Expected: {'sum': 18, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b10011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3241,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 18, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b00001110; cin = 1'b0; // Expected: {'sum': 40, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b00001110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3242,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 40, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b00010110; cin = 1'b1; // Expected: {'sum': 205, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b00010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3243,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 205, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001110; b = 8'b01100110; cin = 1'b1; // Expected: {'sum': 117, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001110; b = 8'b01100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3244,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 117, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010010; b = 8'b00000010; cin = 1'b1; // Expected: {'sum': 85, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010010; b = 8'b00000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3245,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 85, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b01110101; cin = 1'b0; // Expected: {'sum': 225, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b01110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3246,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 225, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b10000101; cin = 1'b0; // Expected: {'sum': 225, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b10000101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3247,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 225, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b11000000; cin = 1'b1; // Expected: {'sum': 133, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b11000000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3248,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 133, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101111; b = 8'b01010110; cin = 1'b0; // Expected: {'sum': 133, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101111; b = 8'b01010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3249,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 133, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b11110111; cin = 1'b0; // Expected: {'sum': 89, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b11110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3250,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 89, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b11000110; cin = 1'b1; // Expected: {'sum': 109, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b11000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3251,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 109, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011010; b = 8'b10011000; cin = 1'b0; // Expected: {'sum': 242, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011010; b = 8'b10011000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3252,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 242, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b11000010; cin = 1'b1; // Expected: {'sum': 48, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b11000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3253,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 48, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b10110011; cin = 1'b0; // Expected: {'sum': 79, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b10110011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3254,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 79, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001000; b = 8'b01111101; cin = 1'b1; // Expected: {'sum': 198, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001000; b = 8'b01111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3255,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 198, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b00011111; cin = 1'b1; // Expected: {'sum': 163, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b00011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3256,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 163, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b11101010; cin = 1'b1; // Expected: {'sum': 5, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b11101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3257,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 5, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b01001100; cin = 1'b1; // Expected: {'sum': 4, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b01001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3258,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b00000010; cin = 1'b0; // Expected: {'sum': 108, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b00000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3259,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 108, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b11011111; cin = 1'b1; // Expected: {'sum': 137, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b11011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3260,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 137, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100111; b = 8'b01011110; cin = 1'b0; // Expected: {'sum': 133, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100111; b = 8'b01011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3261,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 133, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011000; b = 8'b01000001; cin = 1'b0; // Expected: {'sum': 153, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011000; b = 8'b01000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3262,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 153, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100111; b = 8'b10000011; cin = 1'b0; // Expected: {'sum': 234, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100111; b = 8'b10000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3263,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 234, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b00010110; cin = 1'b1; // Expected: {'sum': 81, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b00010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3264,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 81, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b00100110; cin = 1'b1; // Expected: {'sum': 252, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b00100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3265,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 252, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b01010111; cin = 1'b0; // Expected: {'sum': 71, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b01010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3266,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 71, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b10100001; cin = 1'b0; // Expected: {'sum': 3, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b10100001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3267,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001110; b = 8'b01111111; cin = 1'b1; // Expected: {'sum': 142, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001110; b = 8'b01111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3268,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 142, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110101; b = 8'b11010111; cin = 1'b0; // Expected: {'sum': 140, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110101; b = 8'b11010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3269,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 140, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b10000101; cin = 1'b0; // Expected: {'sum': 224, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b10000101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3270,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 224, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b11010010; cin = 1'b0; // Expected: {'sum': 100, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b11010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3271,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 100, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b01011010; cin = 1'b1; // Expected: {'sum': 143, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b01011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3272,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 143, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111000; b = 8'b00100111; cin = 1'b1; // Expected: {'sum': 96, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111000; b = 8'b00100111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3273,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 96, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b11010011; cin = 1'b1; // Expected: {'sum': 42, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b11010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3274,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 42, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b11011011; cin = 1'b1; // Expected: {'sum': 71, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b11011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3275,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 71, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b10000101; cin = 1'b0; // Expected: {'sum': 133, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b10000101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3276,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 133, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b11000010; cin = 1'b1; // Expected: {'sum': 123, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b11000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3277,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 123, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b01101111; cin = 1'b0; // Expected: {'sum': 51, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b01101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3278,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 51, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001000; b = 8'b00101100; cin = 1'b1; // Expected: {'sum': 245, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001000; b = 8'b00101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3279,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 245, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b10011001; cin = 1'b0; // Expected: {'sum': 144, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b10011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3280,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 144, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b11001001; cin = 1'b1; // Expected: {'sum': 124, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b11001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3281,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 124, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101010; b = 8'b11010111; cin = 1'b1; // Expected: {'sum': 130, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101010; b = 8'b11010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3282,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 130, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000100; b = 8'b01000001; cin = 1'b1; // Expected: {'sum': 70, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000100; b = 8'b01000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3283,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 70, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b00001100; cin = 1'b1; // Expected: {'sum': 128, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b00001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3284,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 128, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b11110111; cin = 1'b1; // Expected: {'sum': 28, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b11110111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3285,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 28, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b01111111; cin = 1'b0; // Expected: {'sum': 78, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b01111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3286,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 78, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b10001110; cin = 1'b1; // Expected: {'sum': 229, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b10001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3287,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 229, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b01001001; cin = 1'b0; // Expected: {'sum': 62, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b01001001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3288,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 62, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b10011100; cin = 1'b0; // Expected: {'sum': 116, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b10011100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3289,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 116, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b11110010; cin = 1'b1; // Expected: {'sum': 253, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b11110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3290,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 253, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b10110101; cin = 1'b0; // Expected: {'sum': 225, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b10110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3291,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 225, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100000; b = 8'b01111010; cin = 1'b0; // Expected: {'sum': 154, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100000; b = 8'b01111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3292,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 154, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111011; b = 8'b00100100; cin = 1'b1; // Expected: {'sum': 224, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111011; b = 8'b00100100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3293,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 224, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001111; b = 8'b11010110; cin = 1'b0; // Expected: {'sum': 229, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001111; b = 8'b11010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3294,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 229, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b01011101; cin = 1'b0; // Expected: {'sum': 227, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b01011101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3295,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 227, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010100; b = 8'b10110010; cin = 1'b1; // Expected: {'sum': 135, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010100; b = 8'b10110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3296,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 135, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000111; b = 8'b00100010; cin = 1'b0; // Expected: {'sum': 233, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000111; b = 8'b00100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3297,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 233, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b10110110; cin = 1'b0; // Expected: {'sum': 226, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b10110110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3298,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 226, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b01100000; cin = 1'b1; // Expected: {'sum': 219, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b01100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3299,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 219, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b10001001; cin = 1'b1; // Expected: {'sum': 147, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b10001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3300,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 147, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b01000001; cin = 1'b1; // Expected: {'sum': 252, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b01000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3301,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 252, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b10000101; cin = 1'b1; // Expected: {'sum': 123, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b10000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3302,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 123, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b11000011; cin = 1'b0; // Expected: {'sum': 197, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b11000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3303,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 197, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100001; b = 8'b11100010; cin = 1'b1; // Expected: {'sum': 4, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100001; b = 8'b11100010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3304,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b00111110; cin = 1'b0; // Expected: {'sum': 99, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b00111110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3305,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 99, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111010; b = 8'b10101011; cin = 1'b1; // Expected: {'sum': 166, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111010; b = 8'b10101011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3306,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 166, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100100; b = 8'b10101000; cin = 1'b0; // Expected: {'sum': 76, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100100; b = 8'b10101000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3307,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 76, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011101; b = 8'b00100110; cin = 1'b0; // Expected: {'sum': 3, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011101; b = 8'b00100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3308,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b00010111; cin = 1'b1; // Expected: {'sum': 243, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b00010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3309,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 243, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000100; b = 8'b11100110; cin = 1'b1; // Expected: {'sum': 235, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000100; b = 8'b11100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3310,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 235, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b10010000; cin = 1'b1; // Expected: {'sum': 58, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b10010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3311,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 58, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b10011001; cin = 1'b0; // Expected: {'sum': 230, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b10011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3312,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 230, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b00110010; cin = 1'b0; // Expected: {'sum': 39, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b00110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3313,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 39, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b10110101; cin = 1'b1; // Expected: {'sum': 161, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b10110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3314,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 161, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001000; b = 8'b01100010; cin = 1'b1; // Expected: {'sum': 171, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001000; b = 8'b01100010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3315,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 171, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b11101011; cin = 1'b0; // Expected: {'sum': 189, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b11101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3316,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 189, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001101; b = 8'b11100010; cin = 1'b1; // Expected: {'sum': 240, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001101; b = 8'b11100010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3317,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 240, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b11001010; cin = 1'b1; // Expected: {'sum': 74, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b11001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3318,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 74, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b00110000; cin = 1'b1; // Expected: {'sum': 118, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b00110000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3319,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 118, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b00111111; cin = 1'b0; // Expected: {'sum': 121, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b00111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3320,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 121, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b00101001; cin = 1'b0; // Expected: {'sum': 151, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b00101001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3321,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 151, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b00111010; cin = 1'b0; // Expected: {'sum': 25, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b00111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3322,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 25, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000001; b = 8'b10101010; cin = 1'b0; // Expected: {'sum': 107, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000001; b = 8'b10101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3323,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 107, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b00100101; cin = 1'b0; // Expected: {'sum': 102, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b00100101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3324,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 102, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b01100110; cin = 1'b1; // Expected: {'sum': 64, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b01100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3325,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 64, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b01000110; cin = 1'b1; // Expected: {'sum': 172, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b01000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3326,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 172, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b01111000; cin = 1'b1; // Expected: {'sum': 33, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b01111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3327,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 33, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101001; b = 8'b11001000; cin = 1'b1; // Expected: {'sum': 178, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101001; b = 8'b11001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3328,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 178, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b11100101; cin = 1'b1; // Expected: {'sum': 140, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b11100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3329,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 140, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111111; b = 8'b01111111; cin = 1'b1; // Expected: {'sum': 63, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111111; b = 8'b01111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3330,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 63, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111011; b = 8'b01101111; cin = 1'b0; // Expected: {'sum': 42, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111011; b = 8'b01101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3331,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 42, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b00111101; cin = 1'b0; // Expected: {'sum': 232, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b00111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3332,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 232, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b00111110; cin = 1'b0; // Expected: {'sum': 114, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b00111110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3333,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 114, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011001; b = 8'b00110001; cin = 1'b0; // Expected: {'sum': 138, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011001; b = 8'b00110001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3334,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 138, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001110; b = 8'b01001011; cin = 1'b1; // Expected: {'sum': 154, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001110; b = 8'b01001011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3335,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 154, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b11111101; cin = 1'b1; // Expected: {'sum': 33, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b11111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3336,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 33, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b10010001; cin = 1'b0; // Expected: {'sum': 57, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b10010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3337,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 57, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b10001000; cin = 1'b1; // Expected: {'sum': 218, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b10001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3338,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 218, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101101; b = 8'b01011010; cin = 1'b0; // Expected: {'sum': 7, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101101; b = 8'b01011010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3339,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110111; b = 8'b01010011; cin = 1'b0; // Expected: {'sum': 138, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110111; b = 8'b01010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3340,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 138, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b10010011; cin = 1'b1; // Expected: {'sum': 37, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b10010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3341,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 37, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100000; b = 8'b00011110; cin = 1'b1; // Expected: {'sum': 127, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100000; b = 8'b00011110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3342,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 127, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b10111010; cin = 1'b0; // Expected: {'sum': 244, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b10111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3343,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 244, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b01111101; cin = 1'b1; // Expected: {'sum': 226, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b01111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3344,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 226, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b10011011; cin = 1'b1; // Expected: {'sum': 164, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b10011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3345,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 164, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b11111000; cin = 1'b0; // Expected: {'sum': 157, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b11111000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3346,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 157, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b11100000; cin = 1'b1; // Expected: {'sum': 135, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b11100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3347,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 135, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b10111000; cin = 1'b1; // Expected: {'sum': 221, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b10111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3348,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 221, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b11110111; cin = 1'b0; // Expected: {'sum': 90, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b11110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3349,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 90, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110101; b = 8'b11110100; cin = 1'b1; // Expected: {'sum': 170, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110101; b = 8'b11110100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3350,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 170, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b11101111; cin = 1'b1; // Expected: {'sum': 238, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b11101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3351,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 238, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111011; b = 8'b11110011; cin = 1'b1; // Expected: {'sum': 175, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111011; b = 8'b11110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3352,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 175, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100100; b = 8'b01010011; cin = 1'b1; // Expected: {'sum': 248, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100100; b = 8'b01010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3353,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 248, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110011; b = 8'b01100000; cin = 1'b0; // Expected: {'sum': 19, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110011; b = 8'b01100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3354,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 19, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b01000010; cin = 1'b1; // Expected: {'sum': 46, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b01000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3355,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 46, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b10110111; cin = 1'b0; // Expected: {'sum': 56, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b10110111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3356,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 56, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b01010111; cin = 1'b0; // Expected: {'sum': 132, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b01010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3357,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 132, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b01001111; cin = 1'b0; // Expected: {'sum': 145, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b01001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3358,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 145, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b10001111; cin = 1'b1; // Expected: {'sum': 48, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b10001111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3359,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 48, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b10001001; cin = 1'b1; // Expected: {'sum': 179, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b10001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3360,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 179, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b10001110; cin = 1'b1; // Expected: {'sum': 197, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b10001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3361,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 197, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001101; b = 8'b01001111; cin = 1'b0; // Expected: {'sum': 92, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001101; b = 8'b01001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3362,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 92, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b11011001; cin = 1'b0; // Expected: {'sum': 246, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b11011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3363,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 246, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b01011000; cin = 1'b1; // Expected: {'sum': 141, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b01011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3364,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 141, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b11000000; cin = 1'b0; // Expected: {'sum': 143, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b11000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3365,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 143, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001011; b = 8'b10000111; cin = 1'b1; // Expected: {'sum': 211, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001011; b = 8'b10000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3366,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 211, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b01010000; cin = 1'b1; // Expected: {'sum': 86, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b01010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3367,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 86, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b01000110; cin = 1'b0; // Expected: {'sum': 176, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b01000110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3368,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 176, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101011; b = 8'b11111111; cin = 1'b1; // Expected: {'sum': 43, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101011; b = 8'b11111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3369,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 43, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b00011011; cin = 1'b1; // Expected: {'sum': 64, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b00011011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3370,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 64, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b00101010; cin = 1'b0; // Expected: {'sum': 47, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b00101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3371,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 47, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b10001101; cin = 1'b1; // Expected: {'sum': 149, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b10001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3372,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 149, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b11001101; cin = 1'b1; // Expected: {'sum': 236, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b11001101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3373,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 236, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001000; b = 8'b01111100; cin = 1'b1; // Expected: {'sum': 69, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001000; b = 8'b01111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3374,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 69, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110101; b = 8'b11010001; cin = 1'b1; // Expected: {'sum': 7, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110101; b = 8'b11010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3375,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b10000011; cin = 1'b1; // Expected: {'sum': 208, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b10000011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3376,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 208, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b10100110; cin = 1'b1; // Expected: {'sum': 146, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b10100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3377,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 146, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000110; b = 8'b10000110; cin = 1'b0; // Expected: {'sum': 140, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000110; b = 8'b10000110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3378,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 140, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b10010001; cin = 1'b0; // Expected: {'sum': 108, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b10010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3379,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 108, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001110; b = 8'b11100101; cin = 1'b0; // Expected: {'sum': 51, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001110; b = 8'b11100101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3380,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 51, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b01001111; cin = 1'b1; // Expected: {'sum': 245, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b01001111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3381,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 245, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000101; b = 8'b10100011; cin = 1'b0; // Expected: {'sum': 40, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000101; b = 8'b10100011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3382,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 40, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b11110001; cin = 1'b1; // Expected: {'sum': 163, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b11110001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3383,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 163, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100011; b = 8'b01110111; cin = 1'b1; // Expected: {'sum': 91, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100011; b = 8'b01110111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3384,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 91, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000101; b = 8'b01011111; cin = 1'b0; // Expected: {'sum': 36, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000101; b = 8'b01011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3385,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 36, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000100; b = 8'b10001010; cin = 1'b0; // Expected: {'sum': 142, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000100; b = 8'b10001010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3386,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 142, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000110; b = 8'b11001111; cin = 1'b0; // Expected: {'sum': 21, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000110; b = 8'b11001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3387,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 21, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b01010001; cin = 1'b0; // Expected: {'sum': 82, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b01010001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3388,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 82, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b00100010; cin = 1'b0; // Expected: {'sum': 64, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b00100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3389,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 64, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b00001111; cin = 1'b0; // Expected: {'sum': 247, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b00001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3390,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 247, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101110; b = 8'b11100010; cin = 1'b1; // Expected: {'sum': 17, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101110; b = 8'b11100010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3391,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 17, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b10110110; cin = 1'b1; // Expected: {'sum': 96, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b10110110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3392,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 96, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b01101111; cin = 1'b1; // Expected: {'sum': 241, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b01101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3393,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 241, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b00010111; cin = 1'b0; // Expected: {'sum': 30, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b00010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3394,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 30, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b01010110; cin = 1'b1; // Expected: {'sum': 236, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b01010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3395,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 236, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010101; b = 8'b00110101; cin = 1'b1; // Expected: {'sum': 75, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010101; b = 8'b00110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3396,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 75, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000101; b = 8'b10110010; cin = 1'b0; // Expected: {'sum': 55, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000101; b = 8'b10110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3397,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 55, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b01100000; cin = 1'b0; // Expected: {'sum': 78, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b01100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3398,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 78, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b00100100; cin = 1'b1; // Expected: {'sum': 152, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b00100100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3399,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 152, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b11011100; cin = 1'b0; // Expected: {'sum': 22, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b11011100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3400,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 22, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b10011111; cin = 1'b0; // Expected: {'sum': 159, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b10011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3401,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 159, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111010; b = 8'b01110101; cin = 1'b1; // Expected: {'sum': 112, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111010; b = 8'b01110101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3402,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 112, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b10000011; cin = 1'b0; // Expected: {'sum': 26, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b10000011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3403,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 26, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b10011010; cin = 1'b1; // Expected: {'sum': 60, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b10011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3404,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 60, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b10000011; cin = 1'b1; // Expected: {'sum': 239, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b10000011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3405,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 239, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110001; b = 8'b11111011; cin = 1'b0; // Expected: {'sum': 108, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110001; b = 8'b11111011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3406,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 108, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b01111111; cin = 1'b1; // Expected: {'sum': 64, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b01111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3407,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 64, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b11011000; cin = 1'b1; // Expected: {'sum': 196, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b11011000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3408,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 196, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000100; b = 8'b00001100; cin = 1'b1; // Expected: {'sum': 17, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000100; b = 8'b00001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3409,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 17, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b00101101; cin = 1'b0; // Expected: {'sum': 188, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b00101101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3410,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 188, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b00000101; cin = 1'b1; // Expected: {'sum': 152, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b00000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3411,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 152, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b11100110; cin = 1'b0; // Expected: {'sum': 202, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b11100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3412,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 202, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b10010011; cin = 1'b0; // Expected: {'sum': 133, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b10010011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3413,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 133, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b00010101; cin = 1'b1; // Expected: {'sum': 4, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b00010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3414,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b00010101; cin = 1'b0; // Expected: {'sum': 142, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b00010101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3415,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 142, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b01010101; cin = 1'b1; // Expected: {'sum': 218, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b01010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3416,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 218, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100110; b = 8'b10100010; cin = 1'b1; // Expected: {'sum': 201, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100110; b = 8'b10100010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3417,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 201, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b01110100; cin = 1'b0; // Expected: {'sum': 139, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b01110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3418,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 139, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b00101000; cin = 1'b1; // Expected: {'sum': 63, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b00101000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3419,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 63, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b01100100; cin = 1'b0; // Expected: {'sum': 9, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b01100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3420,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 9, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010010; b = 8'b00111001; cin = 1'b1; // Expected: {'sum': 76, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010010; b = 8'b00111001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3421,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 76, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101001; b = 8'b11101010; cin = 1'b0; // Expected: {'sum': 83, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101001; b = 8'b11101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3422,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 83, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110010; b = 8'b11010101; cin = 1'b0; // Expected: {'sum': 71, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110010; b = 8'b11010101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3423,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 71, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b00010111; cin = 1'b0; // Expected: {'sum': 219, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b00010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3424,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 219, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111110; b = 8'b10001010; cin = 1'b0; // Expected: {'sum': 200, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111110; b = 8'b10001010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3425,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 200, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000011; b = 8'b10101011; cin = 1'b0; // Expected: {'sum': 174, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000011; b = 8'b10101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3426,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 174, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b11101011; cin = 1'b1; // Expected: {'sum': 245, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b11101011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3427,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 245, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101110; b = 8'b00001110; cin = 1'b1; // Expected: {'sum': 189, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101110; b = 8'b00001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3428,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 189, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b01010110; cin = 1'b1; // Expected: {'sum': 96, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b01010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3429,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 96, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100010; b = 8'b01101110; cin = 1'b0; // Expected: {'sum': 16, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100010; b = 8'b01101110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3430,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 16, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b11010100; cin = 1'b1; // Expected: {'sum': 91, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b11010100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3431,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 91, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b11010010; cin = 1'b0; // Expected: {'sum': 61, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b11010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3432,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 61, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b11110001; cin = 1'b0; // Expected: {'sum': 29, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b11110001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3433,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 29, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b00001111; cin = 1'b1; // Expected: {'sum': 60, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b00001111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3434,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 60, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111101; b = 8'b01000010; cin = 1'b0; // Expected: {'sum': 127, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111101; b = 8'b01000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3435,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 127, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b00010001; cin = 1'b1; // Expected: {'sum': 44, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b00010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3436,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 44, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110001; b = 8'b00100001; cin = 1'b1; // Expected: {'sum': 147, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110001; b = 8'b00100001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3437,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 147, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110100; b = 8'b11110101; cin = 1'b0; // Expected: {'sum': 105, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110100; b = 8'b11110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3438,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 105, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001011; b = 8'b01010001; cin = 1'b1; // Expected: {'sum': 157, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001011; b = 8'b01010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3439,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 157, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b10111101; cin = 1'b1; // Expected: {'sum': 141, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b10111101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3440,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 141, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001100; b = 8'b00001100; cin = 1'b1; // Expected: {'sum': 217, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001100; b = 8'b00001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3441,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 217, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b01010100; cin = 1'b1; // Expected: {'sum': 74, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b01010100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3442,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 74, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011111; b = 8'b01000000; cin = 1'b0; // Expected: {'sum': 223, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011111; b = 8'b01000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3443,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 223, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101100; b = 8'b10101101; cin = 1'b0; // Expected: {'sum': 89, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101100; b = 8'b10101101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3444,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 89, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b10100110; cin = 1'b0; // Expected: {'sum': 157, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b10100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3445,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 157, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000001; b = 8'b00011110; cin = 1'b0; // Expected: {'sum': 223, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000001; b = 8'b00011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3446,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 223, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b00001011; cin = 1'b1; // Expected: {'sum': 220, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b00001011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3447,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 220, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000110; b = 8'b01011101; cin = 1'b1; // Expected: {'sum': 100, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000110; b = 8'b01011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3448,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 100, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000110; b = 8'b00111000; cin = 1'b1; // Expected: {'sum': 255, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000110; b = 8'b00111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3449,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 255, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b01010001; cin = 1'b1; // Expected: {'sum': 70, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b01010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3450,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 70, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b11010110; cin = 1'b0; // Expected: {'sum': 175, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b11010110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3451,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 175, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b11111011; cin = 1'b1; // Expected: {'sum': 234, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b11111011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3452,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 234, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b01000110; cin = 1'b1; // Expected: {'sum': 70, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b01000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3453,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 70, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b10111011; cin = 1'b1; // Expected: {'sum': 196, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b10111011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3454,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 196, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b11100001; cin = 1'b0; // Expected: {'sum': 214, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b11100001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3455,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 214, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b11011010; cin = 1'b1; // Expected: {'sum': 255, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b11011010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3456,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 255, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b10001011; cin = 1'b1; // Expected: {'sum': 233, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b10001011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3457,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 233, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b10100001; cin = 1'b0; // Expected: {'sum': 254, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b10100001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3458,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 254, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b00011101; cin = 1'b1; // Expected: {'sum': 37, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b00011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3459,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 37, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b00100111; cin = 1'b1; // Expected: {'sum': 155, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b00100111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3460,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 155, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111101; b = 8'b10100001; cin = 1'b1; // Expected: {'sum': 223, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111101; b = 8'b10100001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3461,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 223, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101111; b = 8'b10101000; cin = 1'b0; // Expected: {'sum': 215, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101111; b = 8'b10101000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3462,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 215, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b11011001; cin = 1'b1; // Expected: {'sum': 122, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b11011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3463,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 122, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011101; b = 8'b00010101; cin = 1'b0; // Expected: {'sum': 242, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011101; b = 8'b00010101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3464,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 242, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b10101000; cin = 1'b0; // Expected: {'sum': 135, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b10101000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3465,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 135, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101111; b = 8'b00110000; cin = 1'b0; // Expected: {'sum': 159, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101111; b = 8'b00110000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3466,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 159, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b10000000; cin = 1'b0; // Expected: {'sum': 255, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b10000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3467,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 255, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110111; b = 8'b11111101; cin = 1'b0; // Expected: {'sum': 52, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110111; b = 8'b11111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3468,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 52, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000101; b = 8'b11111100; cin = 1'b1; // Expected: {'sum': 130, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000101; b = 8'b11111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3469,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 130, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b00111110; cin = 1'b0; // Expected: {'sum': 154, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b00111110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3470,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 154, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b01001111; cin = 1'b0; // Expected: {'sum': 183, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b01001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3471,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 183, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b00011100; cin = 1'b1; // Expected: {'sum': 236, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b00011100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3472,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 236, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b01010100; cin = 1'b0; // Expected: {'sum': 177, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b01010100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3473,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 177, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001100; b = 8'b00101100; cin = 1'b1; // Expected: {'sum': 185, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001100; b = 8'b00101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3474,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 185, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b10110110; cin = 1'b0; // Expected: {'sum': 155, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b10110110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3475,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 155, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010100; b = 8'b10110010; cin = 1'b0; // Expected: {'sum': 134, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010100; b = 8'b10110010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3476,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 134, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b10100000; cin = 1'b0; // Expected: {'sum': 12, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b10100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3477,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001000; b = 8'b00100110; cin = 1'b0; // Expected: {'sum': 238, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001000; b = 8'b00100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3478,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 238, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b10111110; cin = 1'b0; // Expected: {'sum': 242, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b10111110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3479,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 242, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b11011001; cin = 1'b1; // Expected: {'sum': 246, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b11011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3480,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 246, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b10000001; cin = 1'b1; // Expected: {'sum': 228, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b10000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3481,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 228, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b00000110; cin = 1'b1; // Expected: {'sum': 61, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b00000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3482,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 61, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b11110000; cin = 1'b0; // Expected: {'sum': 8, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b11110000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3483,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 8, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101101; b = 8'b11000110; cin = 1'b0; // Expected: {'sum': 115, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101101; b = 8'b11000110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3484,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 115, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b01100011; cin = 1'b1; // Expected: {'sum': 73, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b01100011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3485,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 73, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b01111100; cin = 1'b1; // Expected: {'sum': 205, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b01111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3486,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 205, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b01001001; cin = 1'b0; // Expected: {'sum': 33, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b01001001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3487,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 33, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101111; b = 8'b10111010; cin = 1'b0; // Expected: {'sum': 169, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101111; b = 8'b10111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3488,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 169, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b01100000; cin = 1'b1; // Expected: {'sum': 76, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b01100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3489,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 76, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011111; b = 8'b00001011; cin = 1'b1; // Expected: {'sum': 171, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011111; b = 8'b00001011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3490,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 171, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111101; b = 8'b10101110; cin = 1'b0; // Expected: {'sum': 171, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111101; b = 8'b10101110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3491,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 171, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000101; b = 8'b10010010; cin = 1'b1; // Expected: {'sum': 88, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000101; b = 8'b10010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3492,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 88, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b11001010; cin = 1'b1; // Expected: {'sum': 123, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b11001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3493,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 123, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b10010011; cin = 1'b1; // Expected: {'sum': 48, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b10010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3494,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 48, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010100; b = 8'b11000010; cin = 1'b1; // Expected: {'sum': 151, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010100; b = 8'b11000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3495,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 151, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b10100011; cin = 1'b1; // Expected: {'sum': 7, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b10100011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3496,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b01010101; cin = 1'b1; // Expected: {'sum': 14, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b01010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3497,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001111; b = 8'b10111111; cin = 1'b0; // Expected: {'sum': 206, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001111; b = 8'b10111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3498,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 206, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b11100110; cin = 1'b1; // Expected: {'sum': 9, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b11100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3499,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 9, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111101; b = 8'b00101110; cin = 1'b1; // Expected: {'sum': 44, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111101; b = 8'b00101110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3500,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 44, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011010; b = 8'b00001000; cin = 1'b0; // Expected: {'sum': 98, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011010; b = 8'b00001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3501,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 98, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000000; b = 8'b10101110; cin = 1'b0; // Expected: {'sum': 46, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000000; b = 8'b10101110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3502,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 46, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b01000010; cin = 1'b0; // Expected: {'sum': 235, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b01000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3503,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 235, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001100; b = 8'b10101101; cin = 1'b1; // Expected: {'sum': 186, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001100; b = 8'b10101101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3504,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 186, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100110; b = 8'b00000000; cin = 1'b0; // Expected: {'sum': 102, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100110; b = 8'b00000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3505,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 102, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b10100001; cin = 1'b1; // Expected: {'sum': 30, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b10100001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3506,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 30, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b10001100; cin = 1'b1; // Expected: {'sum': 100, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b10001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3507,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 100, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b10010100; cin = 1'b1; // Expected: {'sum': 249, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b10010100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3508,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 249, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b01111110; cin = 1'b1; // Expected: {'sum': 3, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b01111110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3509,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b01011001; cin = 1'b1; // Expected: {'sum': 24, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b01011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3510,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 24, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100000; b = 8'b10001100; cin = 1'b0; // Expected: {'sum': 172, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100000; b = 8'b10001100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3511,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 172, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000110; b = 8'b00111001; cin = 1'b0; // Expected: {'sum': 255, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000110; b = 8'b00111001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3512,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 255, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b11101101; cin = 1'b0; // Expected: {'sum': 88, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b11101101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3513,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 88, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b00010010; cin = 1'b1; // Expected: {'sum': 213, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b00010010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3514,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 213, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b10011010; cin = 1'b0; // Expected: {'sum': 178, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b10011010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3515,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 178, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000110; b = 8'b00100001; cin = 1'b1; // Expected: {'sum': 40, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000110; b = 8'b00100001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3516,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 40, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100000; b = 8'b01111100; cin = 1'b1; // Expected: {'sum': 157, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100000; b = 8'b01111100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3517,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 157, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b10000010; cin = 1'b0; // Expected: {'sum': 5, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b10000010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3518,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 5, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b11001001; cin = 1'b0; // Expected: {'sum': 37, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b11001001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3519,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 37, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b11110100; cin = 1'b1; // Expected: {'sum': 155, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b11110100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3520,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 155, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110010; b = 8'b01001110; cin = 1'b0; // Expected: {'sum': 192, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110010; b = 8'b01001110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3521,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 192, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011010; b = 8'b11010000; cin = 1'b0; // Expected: {'sum': 170, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011010; b = 8'b11010000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3522,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 170, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b00000000; cin = 1'b0; // Expected: {'sum': 76, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b00000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3523,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 76, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011010; b = 8'b10010011; cin = 1'b1; // Expected: {'sum': 46, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011010; b = 8'b10010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3524,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 46, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b10111011; cin = 1'b1; // Expected: {'sum': 42, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b10111011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3525,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 42, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b11101011; cin = 1'b1; // Expected: {'sum': 74, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b11101011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3526,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 74, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b01010011; cin = 1'b1; // Expected: {'sum': 79, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b01010011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3527,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 79, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100110; b = 8'b11000110; cin = 1'b1; // Expected: {'sum': 45, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100110; b = 8'b11000110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3528,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 45, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b00110110; cin = 1'b0; // Expected: {'sum': 188, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b00110110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3529,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 188, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b11111000; cin = 1'b1; // Expected: {'sum': 17, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b11111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3530,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 17, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001111; b = 8'b10101111; cin = 1'b1; // Expected: {'sum': 191, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001111; b = 8'b10101111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3531,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 191, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b01100111; cin = 1'b1; // Expected: {'sum': 0, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b01100111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3532,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b01111111; cin = 1'b1; // Expected: {'sum': 229, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b01111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3533,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 229, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010010; b = 8'b00101011; cin = 1'b0; // Expected: {'sum': 61, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010010; b = 8'b00101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3534,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 61, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b00011100; cin = 1'b0; // Expected: {'sum': 7, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b00011100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3535,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110111; b = 8'b00000111; cin = 1'b1; // Expected: {'sum': 63, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110111; b = 8'b00000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3536,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 63, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100001; b = 8'b10111011; cin = 1'b1; // Expected: {'sum': 221, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100001; b = 8'b10111011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3537,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 221, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000011; b = 8'b11110010; cin = 1'b1; // Expected: {'sum': 182, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000011; b = 8'b11110010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3538,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 182, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110011; b = 8'b00001000; cin = 1'b1; // Expected: {'sum': 188, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110011; b = 8'b00001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3539,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 188, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b00011001; cin = 1'b1; // Expected: {'sum': 160, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b00011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3540,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 160, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010011; b = 8'b11000000; cin = 1'b1; // Expected: {'sum': 20, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010011; b = 8'b11000000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3541,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 20, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101111; b = 8'b11100110; cin = 1'b0; // Expected: {'sum': 85, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101111; b = 8'b11100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3542,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 85, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b10001100; cin = 1'b0; // Expected: {'sum': 247, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b10001100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3543,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 247, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b01010110; cin = 1'b1; // Expected: {'sum': 2, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b01010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3544,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b10111011; cin = 1'b1; // Expected: {'sum': 173, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b10111011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3545,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 173, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b10000101; cin = 1'b1; // Expected: {'sum': 21, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b10000101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3546,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 21, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101111; b = 8'b01011100; cin = 1'b0; // Expected: {'sum': 139, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101111; b = 8'b01011100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3547,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 139, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b00010101; cin = 1'b1; // Expected: {'sum': 199, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b00010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3548,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 199, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b00101110; cin = 1'b0; // Expected: {'sum': 197, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b00101110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3549,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 197, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010011; b = 8'b11000000; cin = 1'b0; // Expected: {'sum': 147, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010011; b = 8'b11000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3550,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 147, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b11101010; cin = 1'b0; // Expected: {'sum': 123, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b11101010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3551,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 123, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b11011001; cin = 1'b0; // Expected: {'sum': 184, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b11011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3552,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 184, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100000; b = 8'b10100100; cin = 1'b1; // Expected: {'sum': 197, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100000; b = 8'b10100100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3553,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 197, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010100; b = 8'b10010010; cin = 1'b0; // Expected: {'sum': 38, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010100; b = 8'b10010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3554,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 38, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b10110100; cin = 1'b1; // Expected: {'sum': 40, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b10110100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3555,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 40, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b11011110; cin = 1'b0; // Expected: {'sum': 83, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b11011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3556,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 83, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101111; b = 8'b11011111; cin = 1'b0; // Expected: {'sum': 14, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101111; b = 8'b11011111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3557,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101010; b = 8'b11111010; cin = 1'b0; // Expected: {'sum': 164, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101010; b = 8'b11111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3558,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 164, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101001; b = 8'b01001101; cin = 1'b0; // Expected: {'sum': 182, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101001; b = 8'b01001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3559,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 182, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b10011011; cin = 1'b0; // Expected: {'sum': 62, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b10011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3560,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 62, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111011; b = 8'b00110011; cin = 1'b1; // Expected: {'sum': 239, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111011; b = 8'b00110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3561,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 239, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000110; b = 8'b10100110; cin = 1'b1; // Expected: {'sum': 173, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000110; b = 8'b10100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3562,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 173, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100111; b = 8'b10011110; cin = 1'b0; // Expected: {'sum': 133, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100111; b = 8'b10011110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3563,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 133, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101100; b = 8'b10010000; cin = 1'b1; // Expected: {'sum': 61, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101100; b = 8'b10010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3564,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 61, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b01010101; cin = 1'b1; // Expected: {'sum': 140, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b01010101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3565,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 140, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b11010110; cin = 1'b1; // Expected: {'sum': 139, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b11010110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3566,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 139, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b01111000; cin = 1'b0; // Expected: {'sum': 247, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b01111000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3567,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 247, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100110; b = 8'b10001111; cin = 1'b0; // Expected: {'sum': 117, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100110; b = 8'b10001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3568,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 117, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111111; b = 8'b01110000; cin = 1'b1; // Expected: {'sum': 48, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111111; b = 8'b01110000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3569,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 48, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b01010000; cin = 1'b1; // Expected: {'sum': 198, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b01010000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3570,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 198, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110100; b = 8'b01010010; cin = 1'b0; // Expected: {'sum': 198, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110100; b = 8'b01010010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3571,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 198, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b00110110; cin = 1'b0; // Expected: {'sum': 231, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b00110110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3572,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 231, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101110; b = 8'b00101100; cin = 1'b1; // Expected: {'sum': 219, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101110; b = 8'b00101100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3573,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 219, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001000; b = 8'b00011001; cin = 1'b1; // Expected: {'sum': 98, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001000; b = 8'b00011001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3574,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 98, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b01111001; cin = 1'b0; // Expected: {'sum': 152, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b01111001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3575,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 152, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110101; b = 8'b11011011; cin = 1'b0; // Expected: {'sum': 144, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110101; b = 8'b11011011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3576,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 144, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111011; b = 8'b00001000; cin = 1'b1; // Expected: {'sum': 196, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111011; b = 8'b00001000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3577,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 196, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010101; b = 8'b10111110; cin = 1'b0; // Expected: {'sum': 211, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010101; b = 8'b10111110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3578,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 211, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b01000111; cin = 1'b0; // Expected: {'sum': 58, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b01000111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3579,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 58, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b00101110; cin = 1'b1; // Expected: {'sum': 144, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b00101110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3580,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 144, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b10111100; cin = 1'b0; // Expected: {'sum': 61, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b10111100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3581,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 61, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b00110101; cin = 1'b0; // Expected: {'sum': 168, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b00110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3582,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 168, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b10010001; cin = 1'b1; // Expected: {'sum': 27, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b10010001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3583,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 27, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010011; b = 8'b01111011; cin = 1'b1; // Expected: {'sum': 207, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010011; b = 8'b01111011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3584,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 207, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111110; b = 8'b00100000; cin = 1'b1; // Expected: {'sum': 95, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111110; b = 8'b00100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3585,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 95, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100001; b = 8'b01100101; cin = 1'b1; // Expected: {'sum': 135, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100001; b = 8'b01100101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3586,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 135, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b11100101; cin = 1'b0; // Expected: {'sum': 148, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b11100101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3587,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 148, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111111; b = 8'b10011111; cin = 1'b1; // Expected: {'sum': 95, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111111; b = 8'b10011111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3588,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 95, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011001; b = 8'b01000010; cin = 1'b1; // Expected: {'sum': 220, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011001; b = 8'b01000010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3589,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 220, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011010; b = 8'b11001100; cin = 1'b0; // Expected: {'sum': 38, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011010; b = 8'b11001100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3590,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 38, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b11111010; cin = 1'b0; // Expected: {'sum': 16, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b11111010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3591,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 16, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010010; b = 8'b00100000; cin = 1'b0; // Expected: {'sum': 114, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010010; b = 8'b00100000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3592,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 114, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b00111001; cin = 1'b1; // Expected: {'sum': 183, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b00111001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3593,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 183, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000101; b = 8'b01010101; cin = 1'b0; // Expected: {'sum': 26, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000101; b = 8'b01010101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3594,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 26, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b00101111; cin = 1'b0; // Expected: {'sum': 82, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b00101111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3595,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 82, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101001; b = 8'b10101100; cin = 1'b0; // Expected: {'sum': 21, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101001; b = 8'b10101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3596,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 21, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b01101110; cin = 1'b0; // Expected: {'sum': 239, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b01101110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3597,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 239, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b01010111; cin = 1'b1; // Expected: {'sum': 174, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b01010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3598,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 174, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b01100001; cin = 1'b0; // Expected: {'sum': 227, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b01100001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3599,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 227, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100010; b = 8'b01101011; cin = 1'b1; // Expected: {'sum': 14, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100010; b = 8'b01101011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3600,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000111; b = 8'b11000111; cin = 1'b1; // Expected: {'sum': 79, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000111; b = 8'b11000111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3601,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 79, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000111; b = 8'b10011100; cin = 1'b0; // Expected: {'sum': 35, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000111; b = 8'b10011100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3602,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 35, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010010; b = 8'b10001010; cin = 1'b1; // Expected: {'sum': 221, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010010; b = 8'b10001010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3603,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 221, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b01010111; cin = 1'b1; // Expected: {'sum': 138, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b01010111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3604,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 138, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b00000001; cin = 1'b0; // Expected: {'sum': 186, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b00000001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3605,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 186, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111000; b = 8'b11011001; cin = 1'b0; // Expected: {'sum': 209, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111000; b = 8'b11011001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3606,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 209, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110101; b = 8'b11111101; cin = 1'b0; // Expected: {'sum': 178, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110101; b = 8'b11111101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3607,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 178, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b00110011; cin = 1'b1; // Expected: {'sum': 244, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b00110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3608,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 244, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b11100000; cin = 1'b1; // Expected: {'sum': 213, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b11100000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3609,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 213, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001111; b = 8'b11110011; cin = 1'b1; // Expected: {'sum': 67, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001111; b = 8'b11110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3610,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 67, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b11110000; cin = 1'b0; // Expected: {'sum': 225, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b11110000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3611,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 225, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b00110001; cin = 1'b0; // Expected: {'sum': 146, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b00110001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3612,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 146, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110101; b = 8'b11110001; cin = 1'b1; // Expected: {'sum': 39, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110101; b = 8'b11110001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3613,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 39, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b01001000; cin = 1'b0; // Expected: {'sum': 132, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b01001000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3614,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 132, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b01100100; cin = 1'b0; // Expected: {'sum': 51, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b01100100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3615,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 51, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111001; b = 8'b01001111; cin = 1'b0; // Expected: {'sum': 136, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111001; b = 8'b01001111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3616,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 136, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100110; b = 8'b01001101; cin = 1'b0; // Expected: {'sum': 51, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100110; b = 8'b01001101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3617,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 51, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b00100010; cin = 1'b1; // Expected: {'sum': 21, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b00100010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3618,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 21, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b00111110; cin = 1'b0; // Expected: {'sum': 251, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b00111110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3619,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 251, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010100; b = 8'b01000001; cin = 1'b1; // Expected: {'sum': 86, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010100; b = 8'b01000001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3620,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 86, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b10011010; cin = 1'b0; // Expected: {'sum': 145, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b10011010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3621,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 145, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b11100110; cin = 1'b1; // Expected: {'sum': 141, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b11100110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3622,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 141, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b00111110; cin = 1'b1; // Expected: {'sum': 128, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b00111110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3623,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 128, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b10100010; cin = 1'b0; // Expected: {'sum': 108, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b10100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3624,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 108, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b10001111; cin = 1'b1; // Expected: {'sum': 24, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b10001111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3625,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 24, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100111; b = 8'b00001110; cin = 1'b0; // Expected: {'sum': 53, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100111; b = 8'b00001110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3626,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 53, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b10011101; cin = 1'b1; // Expected: {'sum': 127, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b10011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3627,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 127, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b00000101; cin = 1'b0; // Expected: {'sum': 141, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b00000101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3628,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 141, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000011; b = 8'b01001110; cin = 1'b1; // Expected: {'sum': 82, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000011; b = 8'b01001110; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3629,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 82, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b11011101; cin = 1'b1; // Expected: {'sum': 31, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b11011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3630,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 31, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b01101010; cin = 1'b1; // Expected: {'sum': 229, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b01101010; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3631,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 229, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011101; b = 8'b10110100; cin = 1'b0; // Expected: {'sum': 81, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011101; b = 8'b10110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3632,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 81, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011001; b = 8'b10101011; cin = 1'b1; // Expected: {'sum': 69, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011001; b = 8'b10101011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3633,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 69, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b00101100; cin = 1'b0; // Expected: {'sum': 250, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b00101100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3634,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 250, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b01110011; cin = 1'b1; // Expected: {'sum': 140, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b01110011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3635,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 140, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b10111111; cin = 1'b1; // Expected: {'sum': 190, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b10111111; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3636,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 190, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b00111110; cin = 1'b0; // Expected: {'sum': 0, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b00111110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3637,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010101; b = 8'b10101001; cin = 1'b0; // Expected: {'sum': 190, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010101; b = 8'b10101001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3638,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 190, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011010; b = 8'b01111000; cin = 1'b1; // Expected: {'sum': 83, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011010; b = 8'b01111000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3639,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 83, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b10110000; cin = 1'b1; // Expected: {'sum': 199, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b10110000; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3640,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 199, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b11001010; cin = 1'b0; // Expected: {'sum': 10, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b11001010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3641,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b10101001; cin = 1'b0; // Expected: {'sum': 21, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b10101001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3642,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 21, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b00001001; cin = 1'b1; // Expected: {'sum': 87, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b00001001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3643,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 87, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b11101011; cin = 1'b0; // Expected: {'sum': 111, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b11101011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3644,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 111, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b11001100; cin = 1'b1; // Expected: {'sum': 117, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b11001100; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3645,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 117, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b01011101; cin = 1'b1; // Expected: {'sum': 163, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b01011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3646,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 163, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b10010111; cin = 1'b0; // Expected: {'sum': 180, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b10010111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3647,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 180, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b10011101; cin = 1'b1; // Expected: {'sum': 27, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b10011101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3648,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 27, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b01000000; cin = 1'b0; // Expected: {'sum': 140, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b01000000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3649,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 140, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110111; b = 8'b10100110; cin = 1'b0; // Expected: {'sum': 221, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110111; b = 8'b10100110; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3650,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 221, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b01110100; cin = 1'b0; // Expected: {'sum': 12, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b01110100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3651,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101010; b = 8'b00110011; cin = 1'b0; // Expected: {'sum': 29, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101010; b = 8'b00110011; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3652,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 29, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b01100010; cin = 1'b0; // Expected: {'sum': 26, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b01100010; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3653,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 26, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110101; b = 8'b01101101; cin = 1'b1; // Expected: {'sum': 35, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110101; b = 8'b01101101; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3654,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 35, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100111; b = 8'b01111000; cin = 1'b0; // Expected: {'sum': 159, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100111; b = 8'b01111000; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3655,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 159, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011001; b = 8'b01001001; cin = 1'b0; // Expected: {'sum': 226, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011001; b = 8'b01001001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3656,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 226, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b01101001; cin = 1'b1; // Expected: {'sum': 82, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b01101001; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3657,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 82, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b01010100; cin = 1'b0; // Expected: {'sum': 215, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b01010100; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3658,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 215, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b01110101; cin = 1'b0; // Expected: {'sum': 146, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b01110101; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3659,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 146, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b01001001; cin = 1'b0; // Expected: {'sum': 131, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b01001001; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3660,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 131, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b10111111; cin = 1'b0; // Expected: {'sum': 2, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b10111111; cin = 1'b0; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3661,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b11100011; cin = 1'b1; // Expected: {'sum': 143, 'cout': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b11100011; cin = 1'b1; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3662,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 143, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        $finish;
    end
  
endmodule