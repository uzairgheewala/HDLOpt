
`timescale 1ns / 1ps

module tb_N6_adder_subtractor;

    // Parameters
    
    parameter N = 6;
    
     
    // Inputs
    
    reg   cin;
    
    reg  [5:0] i0;
    
    reg  [5:0] i1;
    
    
    // Outputs
    
    wire  [5:0] sum;
    
    
    // Instantiate the Unit Under Test (UUT)
    adder_subtractor  #( N ) uut (
        
        .cin(cin),
        
        .i0(i0),
        
        .i1(i1),
        
        
        .sum(sum)
        
    );

    // Clock generation 
    

    
    
    initial begin
        // Initialize Inputs
        
        cin = 0;
        
        i0 = 0;
        
        i1 = 0;
        
    
        // Wait for global reset
        #100;
    
        // Stimuli
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b101000; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 0,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110111; i1 = 6'b111001; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110111; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 1,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000101; i1 = 6'b101001; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000101; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 2,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b110000; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 3,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b000101; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 4,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000101; i1 = 6'b000000; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000101; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 5,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b001010; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 6,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001000; i1 = 6'b001100; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001000; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 7,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b100011; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 8,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000011; i1 = 6'b000011; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000011; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 9,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101001; i1 = 6'b100111; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101001; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 10,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111000; i1 = 6'b010010; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111000; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 11,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011001; i1 = 6'b000111; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011001; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 12,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b110110; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 13,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100111; i1 = 6'b111101; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100111; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 14,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110011; i1 = 6'b100010; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110011; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 15,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100111; i1 = 6'b100100; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100111; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 16,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b011111; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 17,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b101000; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 18,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b111001; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 19,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000000; i1 = 6'b100000; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000000; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 20,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010100; i1 = 6'b100101; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010100; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 21,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101000; i1 = 6'b101111; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101000; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 22,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000101; i1 = 6'b001011; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000101; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 23,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100110; i1 = 6'b110111; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100110; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 24,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010101; i1 = 6'b110110; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010101; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 25,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b000000; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 26,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b101010; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 27,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001100; i1 = 6'b001001; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001100; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 28,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b100010; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 29,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b010000; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 30,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b101100; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 31,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001110; i1 = 6'b010101; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001110; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 32,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111000; i1 = 6'b111100; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111000; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 33,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b100001; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 34,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010101; i1 = 6'b101110; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010101; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 35,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111100; i1 = 6'b001011; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111100; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 36,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101000; i1 = 6'b111111; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101000; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 37,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010001; i1 = 6'b110111; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010001; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 38,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100100; i1 = 6'b111100; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100100; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 39,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110101; i1 = 6'b011011; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110101; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 40,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000000; i1 = 6'b110101; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000000; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 41,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100100; i1 = 6'b110110; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100100; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 42,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b111111; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 43,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100010; i1 = 6'b110010; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100010; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 44,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101101; i1 = 6'b011110; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101101; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 45,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101011; i1 = 6'b011110; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101011; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 46,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010101; i1 = 6'b110111; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010101; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 47,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b001111; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 48,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010100; i1 = 6'b000001; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010100; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 49,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010000; i1 = 6'b100100; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010000; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 50,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011011; i1 = 6'b100010; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011011; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 51,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b110110; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 52,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b010110; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 53,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101001; i1 = 6'b111000; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101001; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 54,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111010; i1 = 6'b000101; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111010; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 55,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000110; i1 = 6'b110101; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000110; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 56,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001000; i1 = 6'b110110; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001000; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 57,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111110; i1 = 6'b100000; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111110; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 58,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b110100; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 59,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101011; i1 = 6'b011010; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101011; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 60,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001001; i1 = 6'b100011; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001001; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 61,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111111; i1 = 6'b001011; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111111; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 62,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110111; i1 = 6'b111010; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110111; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 63,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010100; i1 = 6'b110110; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010100; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 64,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b110101; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 65,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b101110; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 66,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101011; i1 = 6'b010000; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101011; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 67,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110000; i1 = 6'b010011; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110000; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 68,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100001; i1 = 6'b000011; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100001; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 69,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100110; i1 = 6'b111000; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100110; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 70,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011011; i1 = 6'b010000; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011011; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 71,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b110000; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 72,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b111001; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 73,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010100; i1 = 6'b001101; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010100; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 74,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101101; i1 = 6'b001111; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101101; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 75,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110000; i1 = 6'b110001; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110000; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 76,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b100000; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 77,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000101; i1 = 6'b010000; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000101; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 78,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b010100; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 79,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010001; i1 = 6'b100010; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010001; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 80,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010101; i1 = 6'b011110; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010101; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 81,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111101; i1 = 6'b011111; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111101; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 82,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110001; i1 = 6'b111000; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110001; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 83,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011010; i1 = 6'b101001; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011010; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 84,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011010; i1 = 6'b000100; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011010; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 85,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101101; i1 = 6'b001100; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101101; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 86,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b010001; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 87,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b011010; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 88,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110000; i1 = 6'b000111; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110000; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 89,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100001; i1 = 6'b100101; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100001; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 90,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010000; i1 = 6'b100001; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010000; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 91,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010011; i1 = 6'b101011; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010011; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 92,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000010; i1 = 6'b000010; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000010; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 93,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111111; i1 = 6'b101010; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111111; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 94,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011011; i1 = 6'b111110; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011011; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 95,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101111; i1 = 6'b100111; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101111; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 96,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b010111; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 97,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b111000; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 98,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b001111; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 99,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b100101; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 100,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001110; i1 = 6'b110110; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001110; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 101,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b010111; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 102,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001111; i1 = 6'b010001; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001111; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 103,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b011010; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 104,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010100; i1 = 6'b110010; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010100; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 105,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100001; i1 = 6'b000011; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100001; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 106,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b011110; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 107,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100100; i1 = 6'b000000; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100100; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 108,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b101011; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 109,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011100; i1 = 6'b100111; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011100; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 110,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110001; i1 = 6'b101000; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110001; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 111,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111110; i1 = 6'b001110; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111110; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 112,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100111; i1 = 6'b011011; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100111; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 113,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b101110; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 114,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110000; i1 = 6'b101111; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110000; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 115,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b100100; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 116,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b101000; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 117,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101001; i1 = 6'b000000; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101001; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 118,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b101110; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 119,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010100; i1 = 6'b010000; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010100; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 120,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011010; i1 = 6'b011101; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011010; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 121,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b111100; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 122,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011011; i1 = 6'b000001; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011011; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 123,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111101; i1 = 6'b111010; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111101; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 124,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110001; i1 = 6'b000110; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110001; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 125,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b110110; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 126,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010110; i1 = 6'b011000; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010110; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 127,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000110; i1 = 6'b111000; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000110; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 128,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011110; i1 = 6'b111101; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011110; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 129,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011100; i1 = 6'b001111; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011100; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 130,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111101; i1 = 6'b111001; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111101; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 131,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000101; i1 = 6'b100100; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000101; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 132,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b101011; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 133,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000010; i1 = 6'b001000; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000010; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 134,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101101; i1 = 6'b101001; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101101; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 135,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111010; i1 = 6'b110001; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111010; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 136,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000101; i1 = 6'b111111; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000101; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 137,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001100; i1 = 6'b011101; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001100; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 138,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b010111; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 139,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b010001; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 140,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b011001; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 141,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010101; i1 = 6'b001001; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010101; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 142,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000111; i1 = 6'b100011; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000111; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 143,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111101; i1 = 6'b011101; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111101; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 144,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011000; i1 = 6'b000100; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011000; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 145,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b001011; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 146,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011010; i1 = 6'b001011; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011010; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 147,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010101; i1 = 6'b011101; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010101; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 148,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001110; i1 = 6'b010110; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001110; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 149,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010001; i1 = 6'b001101; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010001; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 150,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001000; i1 = 6'b001011; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001000; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 151,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000010; i1 = 6'b111000; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000010; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 152,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000010; i1 = 6'b000000; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000010; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 153,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010011; i1 = 6'b110101; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010011; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 154,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000110; i1 = 6'b100011; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000110; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 155,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b011110; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 156,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b110110; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 157,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b101001; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 158,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110010; i1 = 6'b110001; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110010; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 159,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101101; i1 = 6'b010111; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101101; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 160,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b011010; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 161,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011111; i1 = 6'b000111; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011111; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 162,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010001; i1 = 6'b010101; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010001; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 163,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011000; i1 = 6'b101011; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011000; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 164,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110111; i1 = 6'b011011; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110111; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 165,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011011; i1 = 6'b010001; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011011; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 166,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110000; i1 = 6'b100001; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110000; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 167,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110100; i1 = 6'b110111; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110100; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 168,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b010111; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 169,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111010; i1 = 6'b110101; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111010; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 170,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110111; i1 = 6'b111100; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110111; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 171,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b111010; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 172,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000110; i1 = 6'b000101; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000110; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 173,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001000; i1 = 6'b100111; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001000; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 174,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b101111; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 175,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010110; i1 = 6'b000111; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010110; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 176,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b010010; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 177,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010100; i1 = 6'b001111; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010100; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 178,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b011100; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 179,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111101; i1 = 6'b110010; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111101; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 180,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110000; i1 = 6'b110011; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110000; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 181,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000111; i1 = 6'b101111; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000111; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 182,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101001; i1 = 6'b101110; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101001; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 183,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101011; i1 = 6'b000010; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101011; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 184,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110100; i1 = 6'b001100; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110100; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 185,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010101; i1 = 6'b001000; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010101; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 186,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110110; i1 = 6'b001011; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110110; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 187,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000100; i1 = 6'b110100; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000100; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 188,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010110; i1 = 6'b010100; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010110; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 189,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111100; i1 = 6'b110001; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111100; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 190,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b000110; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 191,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111110; i1 = 6'b000100; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111110; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 192,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000011; i1 = 6'b101011; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000011; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 193,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010001; i1 = 6'b011010; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010001; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 194,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100100; i1 = 6'b111110; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100100; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 195,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000000; i1 = 6'b011001; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000000; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 196,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b111100; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 197,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b100101; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 198,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101110; i1 = 6'b001000; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101110; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 199,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b101000; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 200,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111010; i1 = 6'b100000; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111010; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 201,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100100; i1 = 6'b111101; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100100; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 202,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010111; i1 = 6'b000111; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010111; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 203,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110001; i1 = 6'b011011; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110001; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 204,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101101; i1 = 6'b111000; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101101; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 205,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101011; i1 = 6'b100100; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101011; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 206,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001000; i1 = 6'b001101; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001000; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 207,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100111; i1 = 6'b001000; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100111; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 208,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b110000; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 209,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b000010; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 210,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010010; i1 = 6'b110100; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010010; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 211,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110101; i1 = 6'b101101; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110101; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 212,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001000; i1 = 6'b011100; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001000; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 213,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011001; i1 = 6'b000100; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011001; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 214,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000000; i1 = 6'b110111; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000000; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 215,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b010010; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 216,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100100; i1 = 6'b110010; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100100; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 217,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110101; i1 = 6'b110100; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110101; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 218,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011100; i1 = 6'b001000; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011100; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 219,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b110101; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 220,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001100; i1 = 6'b010011; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001100; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 221,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010111; i1 = 6'b110001; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010111; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 222,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100001; i1 = 6'b100010; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100001; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 223,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b101001; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 224,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111000; i1 = 6'b101101; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111000; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 225,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b001001; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 226,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101000; i1 = 6'b100100; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101000; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 227,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111010; i1 = 6'b011101; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111010; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 228,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110011; i1 = 6'b101101; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110011; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 229,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b001001; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 230,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b110001; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 231,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b011101; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 232,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b010110; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 233,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b001010; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 234,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b010101; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 235,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001101; i1 = 6'b110110; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001101; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 236,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011011; i1 = 6'b111111; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011011; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 237,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101000; i1 = 6'b000110; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101000; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 238,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111101; i1 = 6'b010111; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111101; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 239,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b011011; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 240,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b010011; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 241,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001110; i1 = 6'b010010; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001110; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 242,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111010; i1 = 6'b011000; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111010; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 243,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b111010; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 244,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b000100; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 245,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011101; i1 = 6'b110010; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011101; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 246,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b000001; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 247,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110101; i1 = 6'b101001; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110101; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 248,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b110110; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 249,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b010101; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 250,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011001; i1 = 6'b111011; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011001; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 251,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000111; i1 = 6'b001011; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000111; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 252,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001100; i1 = 6'b110010; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001100; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 253,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111010; i1 = 6'b010000; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111010; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 254,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000011; i1 = 6'b011110; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000011; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 255,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010011; i1 = 6'b011101; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010011; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 256,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b000001; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 257,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b100111; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 258,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111110; i1 = 6'b011111; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111110; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 259,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b001110; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 260,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b011010; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 261,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110001; i1 = 6'b110010; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110001; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 262,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100100; i1 = 6'b111011; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100100; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 263,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b110010; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 264,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000000; i1 = 6'b000011; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000000; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 265,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000110; i1 = 6'b011001; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000110; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 266,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b001101; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 267,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111101; i1 = 6'b001100; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111101; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 268,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101101; i1 = 6'b000110; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101101; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 269,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b101010; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 270,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b101010; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 271,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b000100; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 272,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001000; i1 = 6'b110001; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001000; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 273,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010101; i1 = 6'b110011; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010101; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 274,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101001; i1 = 6'b011100; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101001; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 275,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110001; i1 = 6'b001011; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110001; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 276,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b001111; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 277,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b100100; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 278,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001100; i1 = 6'b000000; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001100; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 279,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011010; i1 = 6'b000011; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011010; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 280,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b010000; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 281,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110110; i1 = 6'b100010; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110110; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 282,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101011; i1 = 6'b011000; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101011; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 283,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000100; i1 = 6'b001011; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000100; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 284,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111001; i1 = 6'b000011; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111001; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 285,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000110; i1 = 6'b010111; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000110; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 286,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b100100; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 287,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111100; i1 = 6'b001000; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111100; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 288,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111110; i1 = 6'b011100; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111110; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 289,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010110; i1 = 6'b111110; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010110; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 290,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101001; i1 = 6'b111011; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101001; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 291,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b001111; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 292,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110101; i1 = 6'b100000; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110101; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 293,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011101; i1 = 6'b101101; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011101; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 294,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b111000; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 295,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011100; i1 = 6'b111000; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011100; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 296,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010110; i1 = 6'b100000; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010110; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 297,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b000001; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 298,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000000; i1 = 6'b000011; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000000; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 299,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010110; i1 = 6'b100011; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010110; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 300,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111101; i1 = 6'b110011; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111101; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 301,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011011; i1 = 6'b010101; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011011; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 302,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111010; i1 = 6'b100100; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111010; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 303,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001110; i1 = 6'b000100; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001110; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 304,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b111001; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 305,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b010001; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 306,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011011; i1 = 6'b001000; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011011; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 307,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001111; i1 = 6'b000100; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001111; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 308,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b111100; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 309,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101001; i1 = 6'b111100; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101001; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 310,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b110001; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 311,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000111; i1 = 6'b110111; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000111; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 312,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b111011; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 313,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100110; i1 = 6'b101000; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100110; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 314,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101000; i1 = 6'b001111; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101000; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 315,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b100111; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 316,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100001; i1 = 6'b100011; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100001; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 317,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110010; i1 = 6'b000000; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110010; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 318,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b101101; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 319,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110001; i1 = 6'b100100; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110001; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 320,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000000; i1 = 6'b110100; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000000; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 321,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b101010; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 322,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111110; i1 = 6'b001100; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111110; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 323,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b101110; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 324,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011001; i1 = 6'b100000; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011001; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 325,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101111; i1 = 6'b011100; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101111; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 326,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101001; i1 = 6'b111000; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101001; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 327,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b101110; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 328,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111000; i1 = 6'b100011; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111000; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 329,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111001; i1 = 6'b001100; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111001; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 330,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111010; i1 = 6'b110100; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111010; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 331,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111000; i1 = 6'b010101; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111000; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 332,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100011; i1 = 6'b101000; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100011; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 333,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b001101; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 334,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001000; i1 = 6'b000111; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001000; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 335,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b100011; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 336,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001011; i1 = 6'b001110; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001011; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 337,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011111; i1 = 6'b101010; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011111; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 338,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b010100; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 339,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101000; i1 = 6'b111011; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101000; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 340,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b001001; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 341,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b101011; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 342,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011100; i1 = 6'b001101; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011100; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 343,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b000101; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 344,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b010010; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 345,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110011; i1 = 6'b000110; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110011; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 346,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b010000; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 347,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111101; i1 = 6'b100100; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111101; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 348,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101100; i1 = 6'b111010; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101100; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 349,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b110000; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 350,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001011; i1 = 6'b010100; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001011; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 351,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110101; i1 = 6'b000000; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110101; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 352,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000011; i1 = 6'b010100; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000011; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 353,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011001; i1 = 6'b000101; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011001; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 354,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b011111; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 355,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110110; i1 = 6'b000100; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110110; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 356,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101100; i1 = 6'b111111; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101100; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 357,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101110; i1 = 6'b011000; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101110; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 358,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010111; i1 = 6'b111100; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010111; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 359,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111110; i1 = 6'b111011; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111110; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 360,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011000; i1 = 6'b101010; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011000; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 361,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101001; i1 = 6'b000110; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101001; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 362,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011101; i1 = 6'b000100; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011101; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 363,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b000110; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 364,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111000; i1 = 6'b001100; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111000; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 365,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010101; i1 = 6'b001110; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010101; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 366,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001100; i1 = 6'b101111; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001100; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 367,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011000; i1 = 6'b101101; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011000; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 368,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b111110; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 369,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010110; i1 = 6'b000100; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010110; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 370,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101111; i1 = 6'b010111; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101111; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 371,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110110; i1 = 6'b110111; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110110; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 372,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110010; i1 = 6'b111000; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110010; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 373,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b000000; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 374,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111010; i1 = 6'b111101; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111010; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 375,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001111; i1 = 6'b001001; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001111; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 376,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100110; i1 = 6'b001000; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100110; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 377,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101101; i1 = 6'b010101; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101101; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 378,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b001110; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 379,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b010001; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 380,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101110; i1 = 6'b100000; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101110; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 381,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011100; i1 = 6'b110101; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011100; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 382,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101110; i1 = 6'b001111; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101110; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 383,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b110001; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 384,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011100; i1 = 6'b101101; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011100; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 385,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011011; i1 = 6'b110100; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011011; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 386,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001110; i1 = 6'b010001; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001110; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 387,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b010011; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 388,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001000; i1 = 6'b010001; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001000; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 389,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b000101; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 390,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111001; i1 = 6'b101001; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111001; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 391,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110100; i1 = 6'b001000; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110100; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 392,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011001; i1 = 6'b111001; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011001; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 393,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011100; i1 = 6'b010010; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011100; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 394,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000100; i1 = 6'b110010; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000100; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 395,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101110; i1 = 6'b101000; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101110; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 396,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001011; i1 = 6'b010000; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001011; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 397,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001011; i1 = 6'b011010; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001011; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 398,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001100; i1 = 6'b010100; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001100; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 399,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110100; i1 = 6'b101001; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110100; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 400,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001110; i1 = 6'b111001; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001110; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 401,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111100; i1 = 6'b111000; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111100; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 402,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111101; i1 = 6'b101000; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111101; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 403,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011101; i1 = 6'b100110; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011101; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 404,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111111; i1 = 6'b100110; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111111; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 405,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110011; i1 = 6'b110100; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110011; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 406,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101000; i1 = 6'b111001; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101000; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 407,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110111; i1 = 6'b000110; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110111; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 408,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b010001; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 409,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b100110; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 410,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b001010; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 411,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011100; i1 = 6'b110111; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011100; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 412,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010010; i1 = 6'b010010; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010010; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 413,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b011001; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 414,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010101; i1 = 6'b010010; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010101; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 415,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111000; i1 = 6'b011010; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111000; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 416,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111110; i1 = 6'b000001; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111110; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 417,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011110; i1 = 6'b011000; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011110; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 418,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b101101; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 419,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101001; i1 = 6'b110001; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101001; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 420,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010101; i1 = 6'b100010; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010101; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 421,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001101; i1 = 6'b000001; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001101; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 422,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011100; i1 = 6'b100000; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011100; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 423,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010000; i1 = 6'b001100; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010000; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 424,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b111011; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 425,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000011; i1 = 6'b110000; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000011; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 426,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b001101; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 427,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b111101; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 428,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001110; i1 = 6'b010011; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001110; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 429,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100101; i1 = 6'b100001; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100101; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 430,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111100; i1 = 6'b001101; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111100; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 431,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001100; i1 = 6'b111001; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001100; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 432,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b011111; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 433,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010011; i1 = 6'b001001; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010011; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 434,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b110111; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 435,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b111001; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 436,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100011; i1 = 6'b001001; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100011; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 437,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b111000; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 438,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100010; i1 = 6'b110101; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100010; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 439,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010110; i1 = 6'b001011; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010110; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 440,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b001011; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 441,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101011; i1 = 6'b101100; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101011; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 442,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100100; i1 = 6'b000101; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100100; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 443,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111111; i1 = 6'b001110; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111111; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 444,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b110111; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 445,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110010; i1 = 6'b011110; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110010; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 446,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010110; i1 = 6'b110110; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010110; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 447,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b000000; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 448,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001100; i1 = 6'b010101; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001100; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 449,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b010111; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 450,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100100; i1 = 6'b110111; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100100; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 451,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111001; i1 = 6'b001011; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111001; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 452,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110001; i1 = 6'b110100; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110001; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 453,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101001; i1 = 6'b111001; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101001; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 454,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b111101; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 455,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b101000; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 456,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001110; i1 = 6'b000111; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001110; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 457,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b110000; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 458,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011101; i1 = 6'b100100; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011101; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 459,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001000; i1 = 6'b010101; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001000; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 460,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100010; i1 = 6'b011111; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100010; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 461,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b000101; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 462,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100111; i1 = 6'b001100; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100111; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 463,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b101101; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 464,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100001; i1 = 6'b110011; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100001; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 465,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b111011; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 466,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b010001; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 467,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010110; i1 = 6'b100001; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010110; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 468,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111111; i1 = 6'b001000; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111111; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 469,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010101; i1 = 6'b010101; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010101; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 470,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111000; i1 = 6'b111001; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111000; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 471,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011011; i1 = 6'b001001; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011011; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 472,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011111; i1 = 6'b001010; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011111; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 473,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111010; i1 = 6'b101001; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111010; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 474,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100111; i1 = 6'b000000; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100111; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 475,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011011; i1 = 6'b111001; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011011; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 476,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b110111; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 477,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b001111; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 478,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b101100; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 479,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110111; i1 = 6'b111000; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110111; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 480,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010100; i1 = 6'b111001; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010100; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 481,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b111111; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 482,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010110; i1 = 6'b100101; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010110; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 483,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100010; i1 = 6'b011110; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100010; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 484,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100111; i1 = 6'b000111; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100111; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 485,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011010; i1 = 6'b101011; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011010; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 486,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101111; i1 = 6'b100100; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101111; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 487,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101100; i1 = 6'b111001; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101100; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 488,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100101; i1 = 6'b111100; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100101; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 489,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b011101; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 490,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011101; i1 = 6'b111010; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011101; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 491,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111010; i1 = 6'b100110; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111010; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 492,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000010; i1 = 6'b111011; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000010; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 493,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b011101; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 494,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000100; i1 = 6'b000101; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000100; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 495,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011010; i1 = 6'b110111; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011010; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 496,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000011; i1 = 6'b010101; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000011; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 497,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b101011; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 498,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b101110; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 499,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b011011; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 500,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010100; i1 = 6'b011101; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010100; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 501,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110101; i1 = 6'b111111; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110101; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 502,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b101111; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 503,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b101000; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 504,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110100; i1 = 6'b111111; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110100; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 505,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101100; i1 = 6'b001100; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101100; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 506,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111010; i1 = 6'b000101; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111010; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 507,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011101; i1 = 6'b100010; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011101; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 508,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010010; i1 = 6'b010100; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010010; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 509,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110100; i1 = 6'b111110; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110100; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 510,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101101; i1 = 6'b110000; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101101; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 511,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101000; i1 = 6'b101111; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101000; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 512,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000000; i1 = 6'b100001; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000000; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 513,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000101; i1 = 6'b010110; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000101; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 514,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011111; i1 = 6'b100101; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011111; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 515,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111101; i1 = 6'b000010; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111101; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 516,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b110001; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 517,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000111; i1 = 6'b100000; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000111; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 518,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110100; i1 = 6'b111011; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110100; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 519,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b000000; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 520,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b001111; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 521,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011001; i1 = 6'b100100; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011001; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 522,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000110; i1 = 6'b010100; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000110; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 523,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101101; i1 = 6'b011010; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101101; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 524,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000010; i1 = 6'b001111; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000010; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 525,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101110; i1 = 6'b000111; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101110; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 526,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b001110; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 527,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011111; i1 = 6'b111001; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011111; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 528,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000000; i1 = 6'b000110; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000000; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 529,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000000; i1 = 6'b011001; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000000; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 530,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010000; i1 = 6'b000110; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010000; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 531,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101000; i1 = 6'b110100; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101000; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 532,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b001110; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 533,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110000; i1 = 6'b010100; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110000; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 534,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110000; i1 = 6'b110111; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110000; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 535,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011100; i1 = 6'b100010; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011100; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 536,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101101; i1 = 6'b111000; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101101; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 537,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110111; i1 = 6'b011111; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110111; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 538,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010011; i1 = 6'b110111; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010011; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 539,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000000; i1 = 6'b010001; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000000; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 540,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010100; i1 = 6'b010101; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010100; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 541,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010010; i1 = 6'b010111; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010010; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 542,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100101; i1 = 6'b110000; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100101; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 543,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111000; i1 = 6'b010011; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111000; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 544,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010001; i1 = 6'b011000; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010001; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 545,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111010; i1 = 6'b011110; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111010; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 546,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101011; i1 = 6'b111110; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101011; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 547,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b011101; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 548,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100001; i1 = 6'b001001; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100001; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 549,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b111100; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 550,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001011; i1 = 6'b011011; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001011; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 551,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101000; i1 = 6'b001001; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101000; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 552,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110111; i1 = 6'b000101; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110111; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 553,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101100; i1 = 6'b000100; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101100; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 554,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001110; i1 = 6'b000010; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001110; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 555,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b000111; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 556,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010100; i1 = 6'b111111; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010100; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 557,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010001; i1 = 6'b101010; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010001; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 558,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111010; i1 = 6'b000110; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111010; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 559,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011011; i1 = 6'b110100; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011011; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 560,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110101; i1 = 6'b100101; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110101; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 561,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111001; i1 = 6'b000101; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111001; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 562,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110000; i1 = 6'b000110; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110000; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 563,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111110; i1 = 6'b000001; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111110; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 564,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000111; i1 = 6'b000010; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000111; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 565,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110000; i1 = 6'b010000; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110000; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 566,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101111; i1 = 6'b011011; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101111; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 567,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001110; i1 = 6'b110111; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001110; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 568,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b011111; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 569,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b110111; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 570,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b011000; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 571,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b111101; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 572,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000010; i1 = 6'b010101; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000010; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 573,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001111; i1 = 6'b110100; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001111; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 574,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000010; i1 = 6'b010010; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000010; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 575,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100010; i1 = 6'b110000; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100010; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 576,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101011; i1 = 6'b111100; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101011; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 577,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100101; i1 = 6'b110111; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100101; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 578,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b100100; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 579,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b001000; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 580,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011101; i1 = 6'b101010; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011101; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 581,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001110; i1 = 6'b010000; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001110; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 582,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110000; i1 = 6'b001110; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110000; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 583,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111000; i1 = 6'b011001; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111000; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 584,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b011001; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 585,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b000110; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 586,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101011; i1 = 6'b110011; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101011; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 587,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111000; i1 = 6'b001000; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111000; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 588,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101101; i1 = 6'b010001; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101101; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 589,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001000; i1 = 6'b110001; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001000; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 590,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000011; i1 = 6'b001111; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000011; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 591,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011011; i1 = 6'b000101; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011011; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 592,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b110011; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 593,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110111; i1 = 6'b000000; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110111; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 594,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100111; i1 = 6'b000101; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100111; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 595,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111000; i1 = 6'b100110; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111000; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 596,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b011110; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 597,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100110; i1 = 6'b001010; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100110; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 598,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b001100; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 599,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b101111; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 600,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110101; i1 = 6'b011100; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110101; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 601,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b111110; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 602,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101110; i1 = 6'b111100; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101110; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 603,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b110000; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 604,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100101; i1 = 6'b110100; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100101; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 605,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b000010; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 606,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010100; i1 = 6'b011110; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010100; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 607,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110011; i1 = 6'b011101; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110011; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 608,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100100; i1 = 6'b001000; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100100; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 609,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001011; i1 = 6'b101110; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001011; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 610,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b010110; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 611,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111001; i1 = 6'b000111; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111001; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 612,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b011000; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 613,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000110; i1 = 6'b010110; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000110; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 614,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100110; i1 = 6'b111100; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100110; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 615,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010011; i1 = 6'b011001; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010011; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 616,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b101011; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 617,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100001; i1 = 6'b100100; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100001; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 618,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101001; i1 = 6'b000111; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101001; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 619,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000100; i1 = 6'b000110; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000100; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 620,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101101; i1 = 6'b001110; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101101; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 621,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011000; i1 = 6'b100111; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011000; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 622,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001110; i1 = 6'b001101; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001110; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 623,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101011; i1 = 6'b001001; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101011; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 624,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b100000; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 625,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111110; i1 = 6'b100011; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111110; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 626,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100111; i1 = 6'b011011; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100111; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 627,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b011011; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 628,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010111; i1 = 6'b110111; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010111; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 629,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100001; i1 = 6'b011110; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100001; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 630,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b001100; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 631,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100010; i1 = 6'b010100; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100010; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 632,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011110; i1 = 6'b010111; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011110; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 633,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b111111; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 634,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100111; i1 = 6'b001110; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100111; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 635,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100111; i1 = 6'b100111; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100111; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 636,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110110; i1 = 6'b001111; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110110; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 637,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101001; i1 = 6'b011100; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101001; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 638,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b111100; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 639,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b110100; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 640,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b101101; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 641,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010010; i1 = 6'b111001; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010010; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 642,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001001; i1 = 6'b110100; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001001; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 643,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b110010; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 644,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101011; i1 = 6'b100010; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101011; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 645,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011000; i1 = 6'b110101; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011000; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 646,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111010; i1 = 6'b101100; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111010; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 647,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b000110; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 648,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110000; i1 = 6'b001100; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110000; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 649,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110110; i1 = 6'b000010; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110110; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 650,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101001; i1 = 6'b111100; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101001; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 651,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001100; i1 = 6'b001010; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001100; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 652,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001101; i1 = 6'b011010; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001101; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 653,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001110; i1 = 6'b011010; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001110; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 654,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b000111; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 655,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010001; i1 = 6'b110011; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010001; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 656,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101110; i1 = 6'b010100; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101110; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 657,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b011000; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 658,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110011; i1 = 6'b111111; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110011; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 659,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100111; i1 = 6'b001001; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100111; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 660,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b101111; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 661,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000111; i1 = 6'b111000; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000111; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 662,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011011; i1 = 6'b001111; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011011; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 663,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b101101; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 664,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101101; i1 = 6'b100010; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101101; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 665,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b100101; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 666,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001100; i1 = 6'b010101; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001100; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 667,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111000; i1 = 6'b101001; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111000; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 668,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b010111; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 669,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010110; i1 = 6'b111101; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010110; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 670,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101100; i1 = 6'b111000; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101100; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 671,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010101; i1 = 6'b101000; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010101; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 672,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111101; i1 = 6'b000100; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111101; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 673,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110010; i1 = 6'b011010; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110010; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 674,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b011100; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 675,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001100; i1 = 6'b010110; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001100; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 676,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100001; i1 = 6'b111101; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100001; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 677,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101100; i1 = 6'b100101; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101100; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 678,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011101; i1 = 6'b010110; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011101; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 679,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b001100; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 680,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b101001; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 681,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100111; i1 = 6'b000010; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100111; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 682,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110011; i1 = 6'b100011; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110011; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 683,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011110; i1 = 6'b011011; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011110; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 684,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100101; i1 = 6'b011001; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100101; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 685,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011010; i1 = 6'b111010; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011010; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 686,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b110001; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 687,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b001011; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 688,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b110101; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 689,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000110; i1 = 6'b010111; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000110; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 690,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b011011; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 691,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101011; i1 = 6'b111110; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101011; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 692,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100001; i1 = 6'b111111; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100001; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 693,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b101000; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 694,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b100011; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 695,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100001; i1 = 6'b101010; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100001; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 696,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101110; i1 = 6'b001011; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101110; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 697,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000110; i1 = 6'b110110; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000110; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 698,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b000010; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 699,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b000011; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 700,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101110; i1 = 6'b000011; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101110; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 701,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110100; i1 = 6'b010011; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110100; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 702,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110111; i1 = 6'b101010; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110111; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 703,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011010; i1 = 6'b111101; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011010; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 704,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111111; i1 = 6'b000010; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111111; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 705,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000100; i1 = 6'b111000; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000100; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 706,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101111; i1 = 6'b110000; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101111; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 707,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100111; i1 = 6'b011110; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100111; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 708,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101001; i1 = 6'b101101; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101001; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 709,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110011; i1 = 6'b100111; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110011; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 710,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b111111; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 711,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101101; i1 = 6'b011011; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101101; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 712,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001100; i1 = 6'b111000; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001100; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 713,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011001; i1 = 6'b001010; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011001; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 714,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b001101; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 715,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111110; i1 = 6'b110001; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111110; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 716,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111110; i1 = 6'b100110; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111110; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 717,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111010; i1 = 6'b101011; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111010; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 718,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000011; i1 = 6'b010110; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000011; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 719,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100001; i1 = 6'b101111; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100001; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 720,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011100; i1 = 6'b000101; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011100; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 721,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100111; i1 = 6'b001000; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100111; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 722,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b110011; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 723,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000101; i1 = 6'b100010; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000101; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 724,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000110; i1 = 6'b110001; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000110; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 725,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101111; i1 = 6'b101100; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101111; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 726,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100101; i1 = 6'b010111; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100101; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 727,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110010; i1 = 6'b001101; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110010; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 728,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100001; i1 = 6'b010011; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100001; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 729,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101000; i1 = 6'b111001; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101000; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 730,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101000; i1 = 6'b001010; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101000; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 731,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b110010; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 732,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011101; i1 = 6'b011110; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011101; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 733,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110100; i1 = 6'b010011; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110100; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 734,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101110; i1 = 6'b110111; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101110; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 735,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111110; i1 = 6'b000000; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111110; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 736,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101011; i1 = 6'b011101; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101011; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 737,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111110; i1 = 6'b110110; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111110; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 738,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b100110; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 739,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110010; i1 = 6'b001010; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110010; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 740,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011001; i1 = 6'b110101; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011001; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 741,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000111; i1 = 6'b110101; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000111; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 742,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111111; i1 = 6'b111100; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111111; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 743,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011000; i1 = 6'b010100; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011000; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 744,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b111101; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 745,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110011; i1 = 6'b011010; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110011; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 746,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111111; i1 = 6'b111011; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111111; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 747,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111000; i1 = 6'b111000; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111000; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 748,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101101; i1 = 6'b110100; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101101; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 749,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101101; i1 = 6'b001101; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101101; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 750,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000000; i1 = 6'b101010; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000000; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 751,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010001; i1 = 6'b101010; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010001; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 752,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111110; i1 = 6'b011010; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111110; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 753,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b100011; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 754,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101100; i1 = 6'b101110; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101100; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 755,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010111; i1 = 6'b101100; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010111; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 756,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110011; i1 = 6'b111001; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110011; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 757,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001110; i1 = 6'b001101; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001110; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 758,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101100; i1 = 6'b111011; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101100; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 759,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101011; i1 = 6'b001101; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101011; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 760,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011011; i1 = 6'b011111; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011011; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 761,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000000; i1 = 6'b010010; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000000; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 762,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b100000; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 763,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111110; i1 = 6'b000010; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111110; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 764,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110111; i1 = 6'b110000; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110111; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 765,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101001; i1 = 6'b010101; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101001; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 766,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b100100; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 767,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b111110; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 768,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111101; i1 = 6'b100101; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111101; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 769,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111000; i1 = 6'b100100; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111000; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 770,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000110; i1 = 6'b100111; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000110; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 771,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b011110; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 772,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100001; i1 = 6'b000001; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100001; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 773,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b000001; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 774,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b011010; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 775,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111111; i1 = 6'b100110; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111111; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 776,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011001; i1 = 6'b101011; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011001; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 777,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111101; i1 = 6'b010011; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111101; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 778,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111010; i1 = 6'b100100; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111010; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 779,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001110; i1 = 6'b110000; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001110; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 780,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b101000; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 781,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b011000; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 782,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101110; i1 = 6'b110010; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101110; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 783,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101110; i1 = 6'b000100; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101110; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 784,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b001011; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 785,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b001100; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 786,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b101110; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 787,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010100; i1 = 6'b100101; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010100; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 788,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110011; i1 = 6'b101011; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110011; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 789,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000100; i1 = 6'b011000; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000100; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 790,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b101010; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 791,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b000101; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 792,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b110100; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 793,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100011; i1 = 6'b010011; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100011; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 794,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b110001; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 795,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111000; i1 = 6'b000111; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111000; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 796,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100110; i1 = 6'b010111; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100110; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 797,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b000111; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 798,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001111; i1 = 6'b000001; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001111; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 799,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110100; i1 = 6'b011000; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110100; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 800,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101110; i1 = 6'b110100; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101110; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 801,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011001; i1 = 6'b001011; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011001; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 802,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b100100; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 803,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010100; i1 = 6'b010111; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010100; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 804,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111001; i1 = 6'b001101; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111001; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 805,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110011; i1 = 6'b011100; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110011; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 806,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000110; i1 = 6'b111010; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000110; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 807,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b111101; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 808,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b010000; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 809,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011001; i1 = 6'b011101; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011001; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 810,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b101100; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 811,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110110; i1 = 6'b011111; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110110; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 812,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111110; i1 = 6'b010110; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111110; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 813,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000010; i1 = 6'b011010; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000010; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 814,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101011; i1 = 6'b011111; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101011; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 815,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110011; i1 = 6'b001011; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110011; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 816,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100110; i1 = 6'b011111; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100110; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 817,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011011; i1 = 6'b000111; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011011; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 818,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001111; i1 = 6'b101010; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001111; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 819,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011001; i1 = 6'b000010; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011001; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 820,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b010000; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 821,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010011; i1 = 6'b011100; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010011; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 822,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111000; i1 = 6'b100000; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111000; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 823,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101110; i1 = 6'b101000; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101110; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 824,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001000; i1 = 6'b101010; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001000; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 825,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001101; i1 = 6'b010011; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001101; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 826,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111110; i1 = 6'b011111; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111110; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 827,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b110001; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 828,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000100; i1 = 6'b100100; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000100; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 829,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011100; i1 = 6'b011010; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011100; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 830,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b110110; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 831,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100001; i1 = 6'b010001; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100001; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 832,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101101; i1 = 6'b001011; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101101; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 833,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011010; i1 = 6'b000110; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011010; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 834,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010101; i1 = 6'b000000; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010101; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 835,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b010110; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 836,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b001001; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 837,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010101; i1 = 6'b101011; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010101; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 838,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100111; i1 = 6'b111100; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100111; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 839,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011010; i1 = 6'b001001; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011010; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 840,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010010; i1 = 6'b010110; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010010; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 841,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001100; i1 = 6'b011001; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001100; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 842,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010000; i1 = 6'b101110; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010000; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 843,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000110; i1 = 6'b100101; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000110; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 844,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101100; i1 = 6'b100100; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101100; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 845,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b001100; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 846,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110101; i1 = 6'b000100; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110101; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 847,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011001; i1 = 6'b011011; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011001; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 848,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010110; i1 = 6'b101001; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010110; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 849,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111110; i1 = 6'b000110; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111110; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 850,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100010; i1 = 6'b101111; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100010; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 851,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b100000; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 852,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110001; i1 = 6'b100000; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110001; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 853,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b000011; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 854,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b110111; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 855,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000011; i1 = 6'b100111; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000011; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 856,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b100001; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 857,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000000; i1 = 6'b010000; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000000; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 858,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000000; i1 = 6'b001111; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000000; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 859,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000011; i1 = 6'b000111; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000011; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 860,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101011; i1 = 6'b101110; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101011; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 861,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b101011; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 862,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011110; i1 = 6'b010110; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011110; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 863,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000100; i1 = 6'b101001; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000100; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 864,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100001; i1 = 6'b001111; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100001; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 865,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b100001; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 866,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b010011; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 867,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b100101; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 868,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001100; i1 = 6'b011011; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001100; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 869,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b111100; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 870,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011100; i1 = 6'b110010; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011100; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 871,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110010; i1 = 6'b110010; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110010; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 872,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100001; i1 = 6'b101001; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100001; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 873,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b101110; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 874,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110111; i1 = 6'b001111; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110111; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 875,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010010; i1 = 6'b100000; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010010; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 876,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b101011; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 877,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111110; i1 = 6'b000111; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111110; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 878,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b101010; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 879,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b111011; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 880,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110101; i1 = 6'b100001; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110101; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 881,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b101001; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 882,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000110; i1 = 6'b000001; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000110; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 883,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110011; i1 = 6'b111010; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110011; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 884,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011001; i1 = 6'b000001; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011001; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 885,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100101; i1 = 6'b001100; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100101; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 886,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111100; i1 = 6'b010011; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111100; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 887,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b101001; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 888,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b010111; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 889,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b101100; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 890,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110101; i1 = 6'b010000; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110101; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 891,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100111; i1 = 6'b000110; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100111; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 892,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110011; i1 = 6'b100110; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110011; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 893,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011111; i1 = 6'b110110; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011111; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 894,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101111; i1 = 6'b001100; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101111; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 895,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000000; i1 = 6'b001011; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000000; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 896,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110000; i1 = 6'b111100; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110000; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 897,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000111; i1 = 6'b110101; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000111; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 898,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001100; i1 = 6'b000000; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001100; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 899,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b111010; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 900,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b010111; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 901,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011110; i1 = 6'b100110; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011110; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 902,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111101; i1 = 6'b011101; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111101; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 903,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100111; i1 = 6'b001011; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100111; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 904,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110000; i1 = 6'b001000; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110000; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 905,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b010101; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 906,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b110000; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 907,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000111; i1 = 6'b110000; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000111; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 908,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b111001; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 909,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100010; i1 = 6'b011000; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100010; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 910,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111000; i1 = 6'b001111; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111000; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 911,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010111; i1 = 6'b101000; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010111; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 912,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b110011; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 913,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111000; i1 = 6'b010001; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111000; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 914,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b011110; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 915,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010100; i1 = 6'b111110; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010100; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 916,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000000; i1 = 6'b010100; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000000; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 917,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b011011; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 918,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011010; i1 = 6'b110001; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011010; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 919,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b111110; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 920,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011101; i1 = 6'b101000; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011101; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 921,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001100; i1 = 6'b101110; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001100; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 922,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100001; i1 = 6'b011010; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100001; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 923,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010100; i1 = 6'b100001; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010100; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 924,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000000; i1 = 6'b000010; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000000; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 925,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b000100; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 926,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b111101; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 927,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100011; i1 = 6'b010100; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100011; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 928,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100111; i1 = 6'b100011; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100111; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 929,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111110; i1 = 6'b010110; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111110; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 930,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b110000; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 931,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101111; i1 = 6'b101101; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101111; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 932,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b101100; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 933,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b110110; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 934,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110001; i1 = 6'b100110; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110001; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 935,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000111; i1 = 6'b111001; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000111; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 936,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111000; i1 = 6'b100011; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111000; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 937,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b001101; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 938,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b001101; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 939,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100001; i1 = 6'b010000; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100001; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 940,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001000; i1 = 6'b110111; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001000; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 941,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101000; i1 = 6'b001110; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101000; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 942,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101101; i1 = 6'b111011; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101101; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 943,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111110; i1 = 6'b101111; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111110; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 944,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b100101; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 945,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001000; i1 = 6'b100101; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001000; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 946,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110101; i1 = 6'b011000; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110101; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 947,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b001100; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 948,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001100; i1 = 6'b011111; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001100; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 949,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110001; i1 = 6'b000000; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110001; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 950,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011000; i1 = 6'b100000; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011000; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 951,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011101; i1 = 6'b011011; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011101; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 952,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011001; i1 = 6'b101000; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011001; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 953,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010101; i1 = 6'b100110; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010101; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 954,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010100; i1 = 6'b000110; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010100; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 955,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010101; i1 = 6'b001010; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010101; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 956,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000011; i1 = 6'b110010; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000011; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 957,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b110111; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 958,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011011; i1 = 6'b000011; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011011; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 959,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101110; i1 = 6'b000100; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101110; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 960,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b010100; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 961,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000110; i1 = 6'b100001; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000110; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 962,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101001; i1 = 6'b010110; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101001; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 963,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000100; i1 = 6'b110111; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000100; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 964,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010001; i1 = 6'b111000; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010001; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 965,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101101; i1 = 6'b101100; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101101; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 966,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010101; i1 = 6'b011001; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010101; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 967,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111111; i1 = 6'b011110; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111111; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 968,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100001; i1 = 6'b100101; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100001; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 969,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b110111; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 970,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000011; i1 = 6'b110101; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000011; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 971,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b101110; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 972,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b001101; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 973,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001101; i1 = 6'b110100; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001101; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 974,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010110; i1 = 6'b100101; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010110; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 975,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b000101; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 976,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000011; i1 = 6'b110000; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000011; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 977,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001111; i1 = 6'b111001; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001111; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 978,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100111; i1 = 6'b111111; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100111; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 979,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110010; i1 = 6'b110011; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110010; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 980,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b010010; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 981,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b110000; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 982,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001110; i1 = 6'b011100; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001110; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 983,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110011; i1 = 6'b000111; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110011; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 984,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010011; i1 = 6'b110001; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010011; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 985,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110011; i1 = 6'b001111; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110011; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 986,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b100101; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 987,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010100; i1 = 6'b000111; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010100; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 988,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100011; i1 = 6'b111001; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100011; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 989,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100001; i1 = 6'b110100; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100001; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 990,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b110011; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 991,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110100; i1 = 6'b011111; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110100; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 992,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000000; i1 = 6'b000111; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000000; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 993,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001000; i1 = 6'b000001; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001000; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 994,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000101; i1 = 6'b011111; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000101; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 995,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000011; i1 = 6'b000110; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000011; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 996,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110001; i1 = 6'b010101; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110001; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 997,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b001001; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 998,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011001; i1 = 6'b101110; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011001; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 999,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000110; i1 = 6'b001110; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000110; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 1000,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000110; i1 = 6'b001011; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000110; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 1001,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110000; i1 = 6'b101100; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110000; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 1002,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111010; i1 = 6'b101010; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111010; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 1003,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b000010; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 1004,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011001; i1 = 6'b011001; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011001; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 1005,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010110; i1 = 6'b010011; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010110; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 1006,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011011; i1 = 6'b101111; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011011; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 1007,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111100; i1 = 6'b110000; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111100; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 1008,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110011; i1 = 6'b111101; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110011; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 1009,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111100; i1 = 6'b001100; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111100; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 1010,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111010; i1 = 6'b000000; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111010; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 1011,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110001; i1 = 6'b001001; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110001; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 1012,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101101; i1 = 6'b001011; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101101; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 1013,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010100; i1 = 6'b100100; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010100; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 1014,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101000; i1 = 6'b000000; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101000; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 1015,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010010; i1 = 6'b101011; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010010; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 1016,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100100; i1 = 6'b010110; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100100; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 1017,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101000; i1 = 6'b010000; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101000; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 1018,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111111; i1 = 6'b110111; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111111; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 1019,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010110; i1 = 6'b001101; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010110; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 1020,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b000111; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 1021,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111100; i1 = 6'b110100; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111100; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 1022,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110000; i1 = 6'b111000; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110000; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 1023,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010101; i1 = 6'b110100; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010101; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 1024,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b110101; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 1025,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000000; i1 = 6'b111011; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000000; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 1026,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101011; i1 = 6'b000110; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101011; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 1027,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110011; i1 = 6'b000101; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110011; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 1028,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b011010; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 1029,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101001; i1 = 6'b101011; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101001; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 1030,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100111; i1 = 6'b100010; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100111; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 1031,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b100111; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 1032,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111100; i1 = 6'b101110; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111100; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 1033,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110001; i1 = 6'b111110; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110001; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 1034,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b111000; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 1035,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b001001; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 1036,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b111001; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 1037,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010110; i1 = 6'b110101; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010110; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 1038,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b110100; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 1039,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b101100; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 1040,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b100110; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 1041,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101110; i1 = 6'b000111; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101110; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 1042,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011100; i1 = 6'b100001; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011100; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 1043,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b000100; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 1044,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100101; i1 = 6'b001110; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100101; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 1045,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110011; i1 = 6'b110110; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110011; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 1046,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101011; i1 = 6'b100011; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101011; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 1047,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110110; i1 = 6'b100011; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110110; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 1048,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b001011; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 1049,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b001000; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 1050,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101000; i1 = 6'b010100; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101000; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 1051,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110001; i1 = 6'b101110; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110001; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 1052,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b110010; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 1053,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001000; i1 = 6'b000010; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001000; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 1054,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b001010; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 1055,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b001000; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 1056,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111000; i1 = 6'b110011; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111000; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 1057,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011111; i1 = 6'b111101; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011111; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 1058,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011000; i1 = 6'b001100; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011000; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 1059,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000110; i1 = 6'b000000; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000110; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 1060,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b011000; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 1061,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110001; i1 = 6'b111000; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110001; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 1062,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100011; i1 = 6'b010000; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100011; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 1063,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001110; i1 = 6'b101111; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001110; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 1064,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111000; i1 = 6'b100010; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111000; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 1065,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010100; i1 = 6'b111101; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010100; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 1066,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010010; i1 = 6'b100110; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010010; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 1067,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101110; i1 = 6'b101110; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101110; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 1068,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000101; i1 = 6'b100101; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000101; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 1069,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110111; i1 = 6'b011000; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110111; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 1070,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b110100; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 1071,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111010; i1 = 6'b001010; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111010; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 1072,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101011; i1 = 6'b010101; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101011; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 1073,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b000010; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 1074,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001101; i1 = 6'b101101; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001101; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 1075,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000111; i1 = 6'b110110; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000111; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 1076,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b100101; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 1077,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b011010; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 1078,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101100; i1 = 6'b110111; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101100; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 1079,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b101100; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 1080,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010100; i1 = 6'b111000; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010100; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 1081,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b100000; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 1082,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b000010; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 1083,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b111110; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 1084,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101100; i1 = 6'b000100; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101100; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 1085,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001001; i1 = 6'b011001; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001001; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 1086,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b010010; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 1087,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100001; i1 = 6'b100000; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100001; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 1088,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101000; i1 = 6'b111101; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101000; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 1089,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b000010; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 1090,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101001; i1 = 6'b001110; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101001; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 1091,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011111; i1 = 6'b101100; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011111; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 1092,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110000; i1 = 6'b110010; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110000; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 1093,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101100; i1 = 6'b101010; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101100; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 1094,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b010110; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 1095,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010110; i1 = 6'b010011; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010110; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 1096,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b011010; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 1097,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101111; i1 = 6'b000001; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101111; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 1098,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100011; i1 = 6'b000011; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100011; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 1099,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000110; i1 = 6'b001111; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000110; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 1100,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100010; i1 = 6'b000101; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100010; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 1101,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101001; i1 = 6'b010011; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101001; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 1102,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b100000; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 1103,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000110; i1 = 6'b010101; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000110; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 1104,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111111; i1 = 6'b110011; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111111; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 1105,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010010; i1 = 6'b110001; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010010; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 1106,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101011; i1 = 6'b010010; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101011; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 1107,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b001000; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 1108,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010110; i1 = 6'b000001; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010110; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 1109,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101100; i1 = 6'b001101; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101100; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 1110,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001111; i1 = 6'b011110; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001111; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 1111,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110000; i1 = 6'b100000; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110000; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 1112,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b000011; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 1113,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110111; i1 = 6'b000100; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110111; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 1114,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b101000; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 1115,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100001; i1 = 6'b100111; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100001; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 1116,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011011; i1 = 6'b010100; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011011; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 1117,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001100; i1 = 6'b001100; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001100; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 1118,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111111; i1 = 6'b011001; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111111; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 1119,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b100010; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 1120,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110101; i1 = 6'b101111; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110101; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 1121,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101011; i1 = 6'b000010; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101011; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 1122,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000110; i1 = 6'b100100; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000110; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 1123,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b101100; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 1124,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b011010; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 1125,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000111; i1 = 6'b111100; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000111; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 1126,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000000; i1 = 6'b001101; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000000; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 1127,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111000; i1 = 6'b010110; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111000; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 1128,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111110; i1 = 6'b000100; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111110; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 1129,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011001; i1 = 6'b111101; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011001; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 1130,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001001; i1 = 6'b011011; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001001; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 1131,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110111; i1 = 6'b001100; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110111; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 1132,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100001; i1 = 6'b000111; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100001; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 1133,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110001; i1 = 6'b010000; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110001; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 1134,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011001; i1 = 6'b110011; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011001; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 1135,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101110; i1 = 6'b001100; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101110; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 1136,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b010011; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 1137,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b000000; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 1138,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b100001; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 1139,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b101001; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 1140,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111111; i1 = 6'b100010; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111111; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 1141,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001011; i1 = 6'b100101; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001011; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 1142,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100110; i1 = 6'b110001; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100110; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 1143,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010000; i1 = 6'b001111; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010000; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 1144,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000110; i1 = 6'b000110; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000110; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 1145,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000000; i1 = 6'b100110; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000000; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 1146,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101111; i1 = 6'b010011; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101111; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 1147,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101101; i1 = 6'b100000; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101101; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 1148,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011101; i1 = 6'b011111; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011101; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 1149,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111101; i1 = 6'b000010; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111101; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 1150,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b100001; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 1151,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010100; i1 = 6'b101010; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010100; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 1152,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011100; i1 = 6'b101011; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011100; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 1153,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010100; i1 = 6'b001100; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010100; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 1154,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001111; i1 = 6'b011100; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001111; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 1155,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100001; i1 = 6'b100110; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100001; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 1156,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100011; i1 = 6'b111000; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100011; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 1157,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b100001; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 1158,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b101011; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 1159,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000110; i1 = 6'b100010; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000110; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 1160,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010010; i1 = 6'b101101; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010010; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 1161,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001000; i1 = 6'b111011; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001000; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 1162,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b101000; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 1163,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111010; i1 = 6'b111100; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111010; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 1164,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b010010; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 1165,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b011111; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 1166,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010001; i1 = 6'b110100; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010001; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 1167,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110111; i1 = 6'b010100; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110111; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 1168,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010110; i1 = 6'b000010; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010110; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 1169,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010010; i1 = 6'b000111; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010010; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 1170,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011010; i1 = 6'b100010; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011010; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 1171,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b100101; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 1172,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b010100; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 1173,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000000; i1 = 6'b101101; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000000; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 1174,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b101001; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 1175,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111111; i1 = 6'b000010; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111111; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 1176,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100111; i1 = 6'b100001; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100111; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 1177,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101011; i1 = 6'b010110; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101011; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 1178,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111101; i1 = 6'b110101; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111101; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 1179,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b011100; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 1180,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000110; i1 = 6'b001101; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000110; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 1181,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101101; i1 = 6'b001001; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101101; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 1182,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b011111; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 1183,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101100; i1 = 6'b110001; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101100; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 1184,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001011; i1 = 6'b110110; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001011; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 1185,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101000; i1 = 6'b000011; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101000; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 1186,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110010; i1 = 6'b101111; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110010; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 1187,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b110110; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 1188,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b000111; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 1189,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b111111; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 1190,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011101; i1 = 6'b101011; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011101; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 1191,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001100; i1 = 6'b011100; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001100; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 1192,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b011000; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 1193,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111000; i1 = 6'b101011; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111000; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 1194,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000100; i1 = 6'b010011; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000100; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 1195,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111101; i1 = 6'b111101; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111101; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 1196,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111111; i1 = 6'b100011; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111111; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 1197,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b001111; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 1198,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110001; i1 = 6'b001101; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110001; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 1199,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100001; i1 = 6'b011011; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100001; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 1200,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000011; i1 = 6'b001110; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000011; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 1201,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110011; i1 = 6'b110011; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110011; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 1202,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000111; i1 = 6'b011000; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000111; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 1203,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b011001; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 1204,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010010; i1 = 6'b001111; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010010; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 1205,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b011111; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 1206,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011001; i1 = 6'b100110; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011001; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 1207,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110111; i1 = 6'b101111; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110111; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 1208,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101100; i1 = 6'b010011; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101100; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 1209,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110111; i1 = 6'b110100; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110111; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 1210,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b111010; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 1211,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000000; i1 = 6'b100011; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000000; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 1212,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b011011; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 1213,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b111010; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 1214,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100111; i1 = 6'b110010; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100111; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 1215,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101110; i1 = 6'b000110; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101110; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 1216,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101001; i1 = 6'b100001; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101001; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 1217,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101111; i1 = 6'b111011; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101111; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 1218,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111000; i1 = 6'b111011; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111000; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 1219,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111100; i1 = 6'b100110; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111100; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 1220,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110100; i1 = 6'b000100; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110100; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 1221,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b010010; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 1222,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110100; i1 = 6'b110000; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110100; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 1223,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010001; i1 = 6'b111100; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010001; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 1224,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100101; i1 = 6'b010010; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100101; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 1225,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010010; i1 = 6'b001100; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010010; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 1226,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010001; i1 = 6'b110111; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010001; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 1227,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b010001; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 1228,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b011100; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 1229,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110011; i1 = 6'b000100; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110011; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 1230,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101111; i1 = 6'b011001; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101111; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 1231,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011010; i1 = 6'b011110; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011010; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 1232,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b001101; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 1233,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101001; i1 = 6'b110000; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101001; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 1234,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b011010; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 1235,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b001110; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 1236,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000010; i1 = 6'b001010; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000010; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 1237,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101111; i1 = 6'b010010; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101111; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 1238,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b010010; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 1239,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101100; i1 = 6'b111001; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101100; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 1240,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b010111; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 1241,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000110; i1 = 6'b000101; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000110; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 1242,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111101; i1 = 6'b101011; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111101; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 1243,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010100; i1 = 6'b001100; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010100; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 1244,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b001111; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 1245,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b000111; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 1246,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010100; i1 = 6'b011010; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010100; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 1247,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100101; i1 = 6'b110101; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100101; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 1248,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010101; i1 = 6'b101011; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010101; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 1249,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b101101; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 1250,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000011; i1 = 6'b110111; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000011; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 1251,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011101; i1 = 6'b101001; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011101; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 1252,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110111; i1 = 6'b110011; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110111; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 1253,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101011; i1 = 6'b100001; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101011; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 1254,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001000; i1 = 6'b100110; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001000; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 1255,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001101; i1 = 6'b100010; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001101; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 1256,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b100010; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 1257,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000101; i1 = 6'b101010; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000101; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 1258,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b000011; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 1259,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000100; i1 = 6'b010110; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000100; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 1260,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b110011; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 1261,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010101; i1 = 6'b011000; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010101; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 1262,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111100; i1 = 6'b101011; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111100; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 1263,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b010100; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 1264,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110100; i1 = 6'b111101; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110100; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 1265,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001100; i1 = 6'b110110; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001100; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 1266,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001011; i1 = 6'b111001; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001011; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 1267,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101001; i1 = 6'b001111; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101001; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 1268,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010001; i1 = 6'b010100; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010001; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 1269,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110111; i1 = 6'b000001; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110111; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 1270,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b001010; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 1271,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b010110; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 1272,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101000; i1 = 6'b010110; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101000; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 1273,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111010; i1 = 6'b010010; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111010; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 1274,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100100; i1 = 6'b101010; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100100; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 1275,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011011; i1 = 6'b101010; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011011; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 1276,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b001110; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 1277,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100010; i1 = 6'b110100; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100010; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 1278,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111010; i1 = 6'b111010; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111010; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 1279,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000011; i1 = 6'b010101; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000011; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 1280,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b101010; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 1281,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b111000; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 1282,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000011; i1 = 6'b100100; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000011; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 1283,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b100001; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 1284,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011011; i1 = 6'b010001; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011011; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 1285,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b010011; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 1286,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100011; i1 = 6'b100000; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100011; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 1287,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110101; i1 = 6'b111101; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110101; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 1288,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111101; i1 = 6'b100011; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111101; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 1289,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011001; i1 = 6'b001101; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011001; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 1290,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010011; i1 = 6'b001111; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010011; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 1291,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000100; i1 = 6'b001100; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000100; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 1292,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111111; i1 = 6'b111111; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111111; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 1293,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b101100; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 1294,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111101; i1 = 6'b010110; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111101; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 1295,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010011; i1 = 6'b100101; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010011; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 1296,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101001; i1 = 6'b010111; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101001; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 1297,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011000; i1 = 6'b111010; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011000; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 1298,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b100111; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 1299,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b110011; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 1300,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b100100; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 1301,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010101; i1 = 6'b001110; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010101; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 1302,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100010; i1 = 6'b111111; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100010; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 1303,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110001; i1 = 6'b010001; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110001; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 1304,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011111; i1 = 6'b100100; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011111; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 1305,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b001111; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 1306,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b000011; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 1307,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111010; i1 = 6'b010000; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111010; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 1308,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110001; i1 = 6'b100010; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110001; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 1309,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b001101; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 1310,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011010; i1 = 6'b011000; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011010; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 1311,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b000000; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 1312,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100111; i1 = 6'b100100; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100111; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 1313,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101000; i1 = 6'b011010; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101000; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 1314,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111100; i1 = 6'b101000; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111100; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 1315,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b000010; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 1316,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101101; i1 = 6'b011111; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101101; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 1317,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b011101; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 1318,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110000; i1 = 6'b000001; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110000; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 1319,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100111; i1 = 6'b110001; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100111; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 1320,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111010; i1 = 6'b000111; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111010; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 1321,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001100; i1 = 6'b011101; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001100; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 1322,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000011; i1 = 6'b010010; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000011; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 1323,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b100000; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 1324,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001100; i1 = 6'b011010; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001100; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 1325,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101101; i1 = 6'b011001; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101101; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 1326,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111111; i1 = 6'b100100; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111111; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 1327,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111111; i1 = 6'b000110; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111111; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 1328,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101100; i1 = 6'b000110; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101100; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 1329,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011000; i1 = 6'b100010; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011000; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 1330,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110101; i1 = 6'b100101; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110101; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 1331,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010101; i1 = 6'b101010; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010101; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 1332,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111010; i1 = 6'b000010; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111010; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 1333,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000110; i1 = 6'b111101; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000110; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 1334,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b101110; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 1335,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b000001; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 1336,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110011; i1 = 6'b010001; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110011; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 1337,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011010; i1 = 6'b010110; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011010; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 1338,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000011; i1 = 6'b001000; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000011; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 1339,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011011; i1 = 6'b110000; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011011; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 1340,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100111; i1 = 6'b101011; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100111; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 1341,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011111; i1 = 6'b101110; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011111; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 1342,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101000; i1 = 6'b110010; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101000; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 1343,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010000; i1 = 6'b101000; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010000; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 1344,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b000001; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 1345,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b100010; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 1346,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001100; i1 = 6'b000011; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001100; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 1347,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001000; i1 = 6'b001100; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001000; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 1348,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010001; i1 = 6'b011011; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010001; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 1349,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b100111; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 1350,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b001000; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 1351,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b010110; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 1352,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b011101; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 1353,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110000; i1 = 6'b010110; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110000; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 1354,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011100; i1 = 6'b101111; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011100; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 1355,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b101000; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 1356,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101100; i1 = 6'b100100; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101100; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 1357,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b011000; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 1358,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100110; i1 = 6'b101101; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100110; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 1359,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111101; i1 = 6'b101101; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111101; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 1360,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000100; i1 = 6'b010001; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000100; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 1361,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100011; i1 = 6'b000110; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100011; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 1362,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101001; i1 = 6'b110010; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101001; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 1363,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b111000; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 1364,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100100; i1 = 6'b001110; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100100; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 1365,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b000001; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 1366,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000111; i1 = 6'b111011; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000111; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 1367,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011001; i1 = 6'b101111; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011001; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 1368,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010111; i1 = 6'b011011; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010111; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 1369,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101011; i1 = 6'b110001; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101011; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 1370,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010100; i1 = 6'b010110; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010100; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 1371,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110111; i1 = 6'b111011; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110111; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 1372,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b000110; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 1373,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b000011; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 1374,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b111111; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 1375,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b010111; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 1376,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110001; i1 = 6'b110100; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110001; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 1377,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111010; i1 = 6'b101000; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111010; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 1378,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111000; i1 = 6'b110110; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111000; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 1379,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100111; i1 = 6'b100101; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100111; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 1380,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001000; i1 = 6'b100100; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001000; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 1381,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b110100; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 1382,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111110; i1 = 6'b010000; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111110; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 1383,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110010; i1 = 6'b011111; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110010; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 1384,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b010100; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 1385,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000000; i1 = 6'b100100; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000000; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 1386,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111000; i1 = 6'b110001; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111000; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 1387,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100010; i1 = 6'b111010; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100010; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 1388,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111111; i1 = 6'b000011; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111111; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 1389,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b111100; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 1390,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011011; i1 = 6'b111011; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011011; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 1391,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b111101; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 1392,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000111; i1 = 6'b010111; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000111; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 1393,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100110; i1 = 6'b001111; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100110; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 1394,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b101011; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 1395,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110101; i1 = 6'b010100; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110101; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 1396,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101001; i1 = 6'b011101; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101001; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 1397,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101011; i1 = 6'b010011; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101011; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 1398,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b100110; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 1399,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000111; i1 = 6'b111110; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000111; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 1400,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001100; i1 = 6'b110010; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001100; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 1401,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110011; i1 = 6'b001101; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110011; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 1402,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b001111; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 1403,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101110; i1 = 6'b100011; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101110; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 1404,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b111100; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 1405,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111010; i1 = 6'b011111; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111010; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 1406,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000011; i1 = 6'b000110; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000011; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 1407,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101000; i1 = 6'b011101; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101000; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 1408,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b110111; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 1409,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011001; i1 = 6'b011000; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011001; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 1410,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010111; i1 = 6'b001101; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010111; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 1411,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010100; i1 = 6'b010011; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010100; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 1412,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010101; i1 = 6'b110000; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010101; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 1413,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000111; i1 = 6'b000100; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000111; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 1414,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001101; i1 = 6'b001000; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001101; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 1415,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b111001; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 1416,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010000; i1 = 6'b011000; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010000; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 1417,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011000; i1 = 6'b111101; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011000; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 1418,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110000; i1 = 6'b111110; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110000; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 1419,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101011; i1 = 6'b011010; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101011; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 1420,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b001110; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 1421,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101110; i1 = 6'b111010; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101110; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 1422,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b000001; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 1423,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111000; i1 = 6'b000110; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111000; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 1424,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101100; i1 = 6'b001111; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101100; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 1425,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111010; i1 = 6'b110110; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111010; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 1426,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011101; i1 = 6'b010010; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011101; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 1427,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b000000; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 1428,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b000110; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 1429,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b011110; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 1430,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b001011; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 1431,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001001; i1 = 6'b110000; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001001; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 1432,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b000010; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 1433,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010001; i1 = 6'b011111; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010001; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 1434,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010101; i1 = 6'b100001; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010101; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 1435,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101110; i1 = 6'b000000; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101110; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 1436,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110111; i1 = 6'b010011; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110111; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 1437,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110111; i1 = 6'b000101; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110111; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 1438,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b010101; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 1439,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011001; i1 = 6'b011000; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011001; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 1440,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b001111; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 1441,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000100; i1 = 6'b110000; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000100; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 1442,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101011; i1 = 6'b101100; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101011; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 1443,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b111000; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 1444,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100101; i1 = 6'b100100; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100101; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 1445,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000000; i1 = 6'b101101; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000000; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 1446,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b001000; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 1447,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b001100; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 1448,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b111010; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 1449,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001011; i1 = 6'b001001; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001011; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 1450,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011010; i1 = 6'b111101; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011010; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 1451,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b000111; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 1452,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011010; i1 = 6'b000001; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011010; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 1453,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100111; i1 = 6'b001100; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100111; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 1454,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b011010; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 1455,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b010010; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 1456,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b111010; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 1457,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000010; i1 = 6'b111111; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000010; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 1458,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011000; i1 = 6'b100101; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011000; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 1459,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000010; i1 = 6'b111001; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000010; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 1460,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b101100; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 1461,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001000; i1 = 6'b101101; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001000; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 1462,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011110; i1 = 6'b111010; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011110; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 1463,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b111111; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 1464,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100010; i1 = 6'b111100; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100010; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 1465,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110110; i1 = 6'b100111; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110110; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 1466,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100001; i1 = 6'b110110; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100001; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 1467,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001000; i1 = 6'b010100; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001000; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 1468,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110101; i1 = 6'b000101; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110101; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 1469,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001100; i1 = 6'b001110; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001100; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 1470,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b111110; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 1471,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b100101; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 1472,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110101; i1 = 6'b110010; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110101; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 1473,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110100; i1 = 6'b111100; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110100; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 1474,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000011; i1 = 6'b001001; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000011; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 1475,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011001; i1 = 6'b001111; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011001; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 1476,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b010101; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 1477,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b011110; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 1478,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b001001; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 1479,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100010; i1 = 6'b100100; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100010; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 1480,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b111100; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 1481,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111010; i1 = 6'b110001; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111010; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 1482,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111101; i1 = 6'b001001; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111101; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 1483,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111001; i1 = 6'b011101; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111001; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 1484,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011110; i1 = 6'b111011; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011110; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 1485,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100100; i1 = 6'b010001; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100100; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 1486,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101011; i1 = 6'b101110; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101011; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 1487,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000111; i1 = 6'b011010; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000111; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 1488,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001000; i1 = 6'b100111; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001000; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 1489,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010100; i1 = 6'b010100; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010100; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 1490,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001100; i1 = 6'b111000; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001100; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 1491,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110101; i1 = 6'b101000; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110101; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 1492,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011011; i1 = 6'b100001; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011011; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 1493,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b111010; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 1494,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b110110; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 1495,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100100; i1 = 6'b000000; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100100; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 1496,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100010; i1 = 6'b110111; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100010; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 1497,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100111; i1 = 6'b111111; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100111; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 1498,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111001; i1 = 6'b100011; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111001; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 1499,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001101; i1 = 6'b001001; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001101; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 1500,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100010; i1 = 6'b111000; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100010; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 1501,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111111; i1 = 6'b111111; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111111; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 1502,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b011110; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 1503,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010100; i1 = 6'b110100; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010100; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 1504,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110011; i1 = 6'b110001; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110011; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 1505,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100111; i1 = 6'b001010; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100111; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 1506,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111000; i1 = 6'b011101; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111000; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 1507,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b100110; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 1508,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100011; i1 = 6'b100100; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100011; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 1509,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b000100; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 1510,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b000100; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 1511,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b100111; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 1512,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110000; i1 = 6'b001001; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110000; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 1513,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100010; i1 = 6'b100110; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100010; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 1514,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100111; i1 = 6'b001110; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100111; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 1515,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b101101; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 1516,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010000; i1 = 6'b111101; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010000; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 1517,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b011001; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 1518,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b000010; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 1519,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101110; i1 = 6'b100001; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101110; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 1520,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b101101; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 1521,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011001; i1 = 6'b100111; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011001; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 1522,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100101; i1 = 6'b001010; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100101; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 1523,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100110; i1 = 6'b011011; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100110; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 1524,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011100; i1 = 6'b100011; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011100; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 1525,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001011; i1 = 6'b001010; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001011; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 1526,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b001010; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 1527,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101000; i1 = 6'b010111; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101000; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 1528,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011001; i1 = 6'b010000; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011001; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 1529,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b011000; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 1530,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b100110; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 1531,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b100101; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 1532,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100111; i1 = 6'b101101; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100111; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 1533,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b010011; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 1534,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b111011; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 1535,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001100; i1 = 6'b101110; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001100; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 1536,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b011000; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 1537,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001101; i1 = 6'b101111; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001101; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 1538,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000101; i1 = 6'b100011; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000101; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 1539,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000000; i1 = 6'b001010; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000000; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 1540,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100111; i1 = 6'b010010; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100111; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 1541,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110100; i1 = 6'b100011; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110100; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 1542,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010110; i1 = 6'b001101; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010110; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 1543,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b111010; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 1544,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111110; i1 = 6'b001000; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111110; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 1545,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000100; i1 = 6'b001101; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000100; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 1546,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011011; i1 = 6'b001001; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011011; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 1547,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b110110; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 1548,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b110111; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 1549,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111100; i1 = 6'b111111; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111100; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 1550,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b110100; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 1551,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011010; i1 = 6'b100000; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011010; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 1552,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b101010; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 1553,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b110000; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 1554,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b010100; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 1555,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b101011; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 1556,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b000110; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 1557,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010001; i1 = 6'b111111; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010001; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 1558,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011100; i1 = 6'b010011; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011100; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 1559,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101100; i1 = 6'b000000; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101100; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 1560,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011011; i1 = 6'b001011; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011011; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 1561,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111110; i1 = 6'b100100; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111110; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 1562,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111100; i1 = 6'b010110; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111100; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 1563,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b101110; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 1564,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110011; i1 = 6'b111100; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110011; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 1565,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b000100; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 1566,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110100; i1 = 6'b111111; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110100; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 1567,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110100; i1 = 6'b011011; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110100; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 1568,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100100; i1 = 6'b010111; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100100; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 1569,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111111; i1 = 6'b101100; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111111; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 1570,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010001; i1 = 6'b000001; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010001; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 1571,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b011001; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 1572,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000011; i1 = 6'b100001; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000011; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 1573,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101110; i1 = 6'b100101; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101110; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 1574,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110010; i1 = 6'b111101; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110010; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 1575,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010011; i1 = 6'b111110; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010011; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 1576,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000111; i1 = 6'b000011; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000111; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 1577,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110000; i1 = 6'b101110; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110000; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 1578,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011011; i1 = 6'b011011; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011011; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 1579,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011110; i1 = 6'b111100; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011110; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 1580,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101001; i1 = 6'b001001; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101001; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 1581,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011001; i1 = 6'b001101; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011001; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 1582,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b100011; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 1583,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101101; i1 = 6'b100000; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101101; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 1584,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100100; i1 = 6'b111010; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100100; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 1585,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b110011; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 1586,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b000011; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 1587,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110001; i1 = 6'b011111; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110001; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 1588,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b001010; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 1589,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011001; i1 = 6'b011111; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011001; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 1590,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000101; i1 = 6'b111100; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000101; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 1591,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b001100; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 1592,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100101; i1 = 6'b001001; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100101; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 1593,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b000101; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 1594,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b100101; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 1595,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101101; i1 = 6'b111001; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101101; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 1596,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101100; i1 = 6'b100001; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101100; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 1597,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b100000; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 1598,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b111000; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 1599,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111101; i1 = 6'b110110; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111101; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 1600,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b100010; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 1601,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110101; i1 = 6'b101100; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110101; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 1602,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010111; i1 = 6'b000000; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010111; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 1603,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010100; i1 = 6'b011000; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010100; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 1604,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110001; i1 = 6'b000000; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110001; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 1605,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b101111; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 1606,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110111; i1 = 6'b011101; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110111; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 1607,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101001; i1 = 6'b111111; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101001; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 1608,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010111; i1 = 6'b101010; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010111; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 1609,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110111; i1 = 6'b100000; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110111; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 1610,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100001; i1 = 6'b111011; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100001; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 1611,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b110110; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 1612,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110100; i1 = 6'b001010; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110100; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 1613,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101100; i1 = 6'b100110; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101100; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 1614,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101110; i1 = 6'b000001; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101110; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 1615,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011101; i1 = 6'b000111; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011101; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 1616,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000100; i1 = 6'b111111; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000100; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 1617,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000100; i1 = 6'b010111; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000100; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 1618,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111100; i1 = 6'b000001; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111100; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 1619,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010000; i1 = 6'b110001; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010000; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 1620,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110001; i1 = 6'b001010; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110001; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 1621,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111000; i1 = 6'b110101; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111000; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 1622,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110101; i1 = 6'b110110; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110101; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 1623,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001011; i1 = 6'b110111; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001011; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 1624,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001000; i1 = 6'b101000; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001000; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 1625,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100001; i1 = 6'b011111; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100001; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 1626,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101011; i1 = 6'b111011; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101011; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 1627,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b001100; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 1628,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b110101; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 1629,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b110010; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 1630,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110111; i1 = 6'b101110; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110111; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 1631,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b010110; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 1632,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000100; i1 = 6'b110001; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000100; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 1633,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110101; i1 = 6'b010101; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110101; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 1634,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111100; i1 = 6'b111100; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111100; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 1635,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001001; i1 = 6'b010110; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001001; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 1636,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010100; i1 = 6'b100110; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010100; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 1637,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b110101; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 1638,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000000; i1 = 6'b001011; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000000; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 1639,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b100011; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 1640,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010101; i1 = 6'b101000; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010101; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 1641,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111001; i1 = 6'b001001; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111001; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 1642,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010111; i1 = 6'b010000; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010111; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 1643,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011100; i1 = 6'b000000; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011100; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 1644,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010110; i1 = 6'b100010; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010110; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 1645,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b010000; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 1646,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111010; i1 = 6'b001110; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111010; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 1647,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001011; i1 = 6'b001000; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001011; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 1648,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101001; i1 = 6'b001001; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101001; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 1649,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110011; i1 = 6'b010110; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110011; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 1650,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010110; i1 = 6'b010110; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010110; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 1651,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b100011; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 1652,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b011011; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 1653,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b011100; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 1654,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000100; i1 = 6'b110101; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000100; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 1655,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b101111; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 1656,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000000; i1 = 6'b111011; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000000; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 1657,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b011110; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 1658,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110010; i1 = 6'b111100; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110010; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 1659,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110001; i1 = 6'b100000; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110001; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 1660,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b110100; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 1661,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b010000; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 1662,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001100; i1 = 6'b010110; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001100; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 1663,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b001010; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 1664,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110011; i1 = 6'b100110; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110011; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 1665,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101100; i1 = 6'b100001; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101100; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 1666,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001110; i1 = 6'b110111; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001110; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 1667,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b100011; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 1668,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b001011; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 1669,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b101011; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 1670,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100010; i1 = 6'b100000; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100010; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 1671,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b001010; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 1672,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110111; i1 = 6'b001001; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110111; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 1673,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011100; i1 = 6'b010011; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011100; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 1674,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b110000; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 1675,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b001001; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 1676,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b100110; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 1677,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101110; i1 = 6'b000011; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101110; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 1678,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b110011; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 1679,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011001; i1 = 6'b111110; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011001; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 1680,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111100; i1 = 6'b101010; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111100; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 1681,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000000; i1 = 6'b110011; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000000; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 1682,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000100; i1 = 6'b011010; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000100; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 1683,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110110; i1 = 6'b111111; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110110; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 1684,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010000; i1 = 6'b011111; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010000; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 1685,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101000; i1 = 6'b010001; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101000; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 1686,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b010100; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 1687,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111010; i1 = 6'b010110; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111010; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 1688,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b010001; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 1689,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010001; i1 = 6'b100011; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010001; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 1690,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b010100; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 1691,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b100101; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 1692,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011000; i1 = 6'b101000; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011000; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 1693,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100011; i1 = 6'b110101; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100011; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 1694,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b100010; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 1695,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110111; i1 = 6'b101100; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110111; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 1696,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111100; i1 = 6'b000111; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111100; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 1697,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100100; i1 = 6'b001111; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100100; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 1698,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100001; i1 = 6'b110000; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100001; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 1699,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100100; i1 = 6'b000111; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100100; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 1700,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001000; i1 = 6'b010110; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001000; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 1701,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100100; i1 = 6'b001100; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100100; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 1702,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011001; i1 = 6'b010010; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011001; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 1703,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b110010; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 1704,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100111; i1 = 6'b110000; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100111; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 1705,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b110011; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 1706,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000010; i1 = 6'b110010; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000010; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 1707,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111010; i1 = 6'b011000; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111010; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 1708,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000111; i1 = 6'b101101; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000111; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 1709,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b010011; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 1710,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b111111; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 1711,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001111; i1 = 6'b101100; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001111; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 1712,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001000; i1 = 6'b110101; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001000; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 1713,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b000100; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 1714,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100010; i1 = 6'b110001; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100010; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 1715,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b000011; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 1716,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b011101; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 1717,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b110010; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 1718,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110000; i1 = 6'b111000; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110000; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 1719,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b001010; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 1720,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010010; i1 = 6'b000101; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010010; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 1721,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011001; i1 = 6'b011110; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011001; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 1722,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001001; i1 = 6'b100000; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001001; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 1723,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111111; i1 = 6'b011100; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111111; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 1724,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011010; i1 = 6'b010110; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011010; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 1725,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b000101; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 1726,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100010; i1 = 6'b101111; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100010; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 1727,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100100; i1 = 6'b010100; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100100; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 1728,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001111; i1 = 6'b110001; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001111; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 1729,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111000; i1 = 6'b100111; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111000; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 1730,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000100; i1 = 6'b010100; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000100; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 1731,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111001; i1 = 6'b010110; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111001; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 1732,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b000000; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 1733,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100010; i1 = 6'b011110; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100010; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 1734,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b010101; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 1735,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001100; i1 = 6'b110011; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001100; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 1736,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000111; i1 = 6'b110001; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000111; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 1737,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000000; i1 = 6'b111010; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000000; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 1738,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111111; i1 = 6'b001000; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111111; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 1739,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b111100; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 1740,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010101; i1 = 6'b111101; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010101; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 1741,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b001100; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 1742,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110111; i1 = 6'b000111; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110111; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 1743,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b100001; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 1744,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111110; i1 = 6'b101011; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111110; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 1745,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110110; i1 = 6'b100101; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110110; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 1746,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011101; i1 = 6'b101001; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011101; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 1747,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011000; i1 = 6'b110010; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011000; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 1748,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110100; i1 = 6'b011001; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110100; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 1749,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001111; i1 = 6'b010110; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001111; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 1750,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101100; i1 = 6'b101100; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101100; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 1751,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101111; i1 = 6'b111001; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101111; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 1752,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b110010; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 1753,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b010010; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 1754,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111101; i1 = 6'b001101; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111101; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 1755,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b001011; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 1756,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111010; i1 = 6'b001111; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111010; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 1757,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100100; i1 = 6'b111010; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100100; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 1758,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111000; i1 = 6'b100100; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111000; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 1759,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010001; i1 = 6'b111000; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010001; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 1760,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011111; i1 = 6'b110111; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011111; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 1761,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001110; i1 = 6'b001010; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001110; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 1762,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b101111; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 1763,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b011001; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 1764,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111010; i1 = 6'b111001; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111010; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 1765,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100110; i1 = 6'b010011; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100110; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 1766,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000111; i1 = 6'b111010; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000111; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 1767,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111000; i1 = 6'b111101; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111000; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 1768,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011101; i1 = 6'b001010; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011101; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 1769,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b111010; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 1770,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b000001; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 1771,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011110; i1 = 6'b101100; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011110; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 1772,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010011; i1 = 6'b011000; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010011; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 1773,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b010111; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 1774,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111101; i1 = 6'b110000; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111101; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 1775,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000000; i1 = 6'b111101; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000000; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 1776,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001100; i1 = 6'b100100; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001100; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 1777,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b010110; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 1778,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111010; i1 = 6'b101110; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111010; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 1779,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b101100; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 1780,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010111; i1 = 6'b101111; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010111; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 1781,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010111; i1 = 6'b000110; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010111; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 1782,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010101; i1 = 6'b101100; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010101; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 1783,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001110; i1 = 6'b010000; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001110; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 1784,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000101; i1 = 6'b110011; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000101; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 1785,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b000110; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 1786,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111111; i1 = 6'b010100; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111111; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 1787,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b110001; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 1788,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111001; i1 = 6'b010100; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111001; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 1789,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011101; i1 = 6'b000111; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011101; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 1790,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100010; i1 = 6'b011010; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100010; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 1791,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011111; i1 = 6'b011100; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011111; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 1792,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111111; i1 = 6'b000100; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111111; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 1793,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b111010; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 1794,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b000011; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 1795,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000110; i1 = 6'b100000; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000110; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 1796,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110010; i1 = 6'b001110; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110010; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 1797,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111111; i1 = 6'b010110; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111111; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 1798,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011001; i1 = 6'b011010; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011001; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 1799,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011000; i1 = 6'b001011; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011000; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 1800,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001110; i1 = 6'b101010; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001110; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 1801,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110000; i1 = 6'b001111; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110000; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 1802,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b111010; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 1803,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b010001; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 1804,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b101111; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 1805,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b011111; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 1806,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101011; i1 = 6'b001000; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101011; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 1807,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010100; i1 = 6'b011111; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010100; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 1808,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b001010; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 1809,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110101; i1 = 6'b001000; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110101; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 1810,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110110; i1 = 6'b111101; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110110; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 1811,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101011; i1 = 6'b101111; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101011; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 1812,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111010; i1 = 6'b001101; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111010; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 1813,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b010011; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 1814,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011101; i1 = 6'b010111; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011101; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 1815,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b101001; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 1816,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101101; i1 = 6'b011101; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101101; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 1817,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b001111; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 1818,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b110001; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 1819,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101101; i1 = 6'b001101; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101101; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 1820,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b110100; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 1821,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b000010; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 1822,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b110011; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 1823,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110001; i1 = 6'b101011; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110001; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 1824,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001100; i1 = 6'b010011; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001100; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 1825,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b010111; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 1826,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100111; i1 = 6'b111101; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100111; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 1827,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b101001; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 1828,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110110; i1 = 6'b111011; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110110; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 1829,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b000010; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 1830,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010001; i1 = 6'b010000; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010001; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 1831,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010001; i1 = 6'b100111; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010001; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 1832,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011110; i1 = 6'b110111; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011110; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 1833,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b110100; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 1834,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000000; i1 = 6'b101111; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000000; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 1835,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001101; i1 = 6'b000101; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001101; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 1836,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100010; i1 = 6'b001101; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100010; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 1837,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101001; i1 = 6'b000111; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101001; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 1838,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b011010; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 1839,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011011; i1 = 6'b100000; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011011; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 1840,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001011; i1 = 6'b110100; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001011; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 1841,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011111; i1 = 6'b110010; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011111; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 1842,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010001; i1 = 6'b110000; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010001; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 1843,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b001110; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 1844,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100011; i1 = 6'b101110; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100011; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 1845,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b100110; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 1846,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001001; i1 = 6'b110010; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001001; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 1847,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000010; i1 = 6'b100101; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000010; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 1848,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010001; i1 = 6'b100001; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010001; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 1849,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110101; i1 = 6'b101110; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110101; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 1850,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010001; i1 = 6'b110100; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010001; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 1851,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b011011; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 1852,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000010; i1 = 6'b000001; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000010; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 1853,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b100100; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 1854,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b101100; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 1855,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b011010; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 1856,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100111; i1 = 6'b011000; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100111; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 1857,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000000; i1 = 6'b001111; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000000; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 1858,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100111; i1 = 6'b011100; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100111; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 1859,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111000; i1 = 6'b000011; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111000; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 1860,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100101; i1 = 6'b010011; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100101; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 1861,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110111; i1 = 6'b101011; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110111; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 1862,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b011001; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 1863,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101001; i1 = 6'b110111; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101001; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 1864,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001101; i1 = 6'b010100; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001101; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 1865,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011011; i1 = 6'b100011; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011011; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 1866,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011110; i1 = 6'b001001; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011110; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 1867,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101000; i1 = 6'b100000; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101000; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 1868,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b101010; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 1869,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111100; i1 = 6'b100100; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111100; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 1870,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010001; i1 = 6'b100110; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010001; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 1871,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111111; i1 = 6'b000011; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111111; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 1872,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b111111; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 1873,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111001; i1 = 6'b110101; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111001; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 1874,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001111; i1 = 6'b001010; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001111; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 1875,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011101; i1 = 6'b011101; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011101; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 1876,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010011; i1 = 6'b010110; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010011; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 1877,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111110; i1 = 6'b011011; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111110; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 1878,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b100111; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 1879,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b101100; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 1880,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b011010; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 1881,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010010; i1 = 6'b101100; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010010; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 1882,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b111010; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 1883,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110111; i1 = 6'b111001; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110111; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 1884,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b111010; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 1885,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b010010; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 1886,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000110; i1 = 6'b001001; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000110; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 1887,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b101101; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 1888,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100001; i1 = 6'b011000; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100001; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 1889,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b011011; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 1890,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b101010; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 1891,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001110; i1 = 6'b100110; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001110; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 1892,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b001111; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 1893,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b101100; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 1894,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111110; i1 = 6'b010001; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111110; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 1895,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011011; i1 = 6'b001010; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011011; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 1896,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001110; i1 = 6'b110100; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001110; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 1897,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010110; i1 = 6'b110000; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010110; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 1898,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000111; i1 = 6'b100000; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000111; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 1899,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b101101; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 1900,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100011; i1 = 6'b100001; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100011; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 1901,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110001; i1 = 6'b110101; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110001; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 1902,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b111010; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 1903,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100100; i1 = 6'b011000; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100100; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 1904,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001000; i1 = 6'b111100; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001000; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 1905,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111111; i1 = 6'b101100; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111111; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 1906,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001111; i1 = 6'b001011; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001111; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 1907,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110110; i1 = 6'b010010; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110110; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 1908,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100011; i1 = 6'b110000; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100011; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 1909,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000111; i1 = 6'b111111; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000111; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 1910,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b110100; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 1911,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b001100; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 1912,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101000; i1 = 6'b111000; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101000; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 1913,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110111; i1 = 6'b101000; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110111; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 1914,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b000100; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 1915,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b101100; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 1916,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b001000; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 1917,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101110; i1 = 6'b101010; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101110; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 1918,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101000; i1 = 6'b110011; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101000; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 1919,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b100111; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 1920,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111101; i1 = 6'b100111; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111101; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 1921,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001011; i1 = 6'b000101; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001011; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 1922,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110000; i1 = 6'b000100; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110000; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 1923,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010011; i1 = 6'b110000; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010011; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 1924,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b110100; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 1925,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000011; i1 = 6'b100010; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000011; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 1926,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b011001; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 1927,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b011011; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 1928,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011111; i1 = 6'b001101; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011111; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 1929,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111001; i1 = 6'b011110; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111001; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 1930,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011110; i1 = 6'b000111; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011110; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 1931,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011001; i1 = 6'b000011; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011001; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 1932,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101100; i1 = 6'b100101; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101100; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 1933,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111010; i1 = 6'b011111; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111010; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 1934,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101001; i1 = 6'b101001; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101001; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 1935,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101100; i1 = 6'b001010; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101100; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 1936,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b111110; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 1937,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110101; i1 = 6'b111101; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110101; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 1938,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b101111; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 1939,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011000; i1 = 6'b000010; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011000; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 1940,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b011010; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 1941,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010010; i1 = 6'b100100; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010010; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 1942,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010001; i1 = 6'b100101; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010001; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 1943,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101100; i1 = 6'b001001; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101100; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 1944,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000000; i1 = 6'b010111; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000000; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 1945,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001011; i1 = 6'b111011; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001011; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 1946,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b101001; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 1947,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100001; i1 = 6'b001100; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100001; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 1948,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100001; i1 = 6'b001010; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100001; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 1949,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001100; i1 = 6'b000100; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001100; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 1950,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b100111; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 1951,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b011110; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 1952,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b101111; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 1953,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101000; i1 = 6'b101101; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101000; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 1954,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b010011; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 1955,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111111; i1 = 6'b000001; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111111; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 1956,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001101; i1 = 6'b101010; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001101; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 1957,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011100; i1 = 6'b000001; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011100; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 1958,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101101; i1 = 6'b010111; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101101; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 1959,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b100100; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 1960,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011101; i1 = 6'b111011; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011101; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 1961,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101110; i1 = 6'b000101; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101110; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 1962,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b011011; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 1963,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000011; i1 = 6'b101100; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000011; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 1964,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b001110; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 1965,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010001; i1 = 6'b111001; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010001; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 1966,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b010000; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 1967,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101111; i1 = 6'b000000; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101111; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 1968,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b101011; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 1969,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011110; i1 = 6'b100000; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011110; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 1970,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100110; i1 = 6'b000100; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100110; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 1971,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011001; i1 = 6'b110100; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011001; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 1972,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b000101; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 1973,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b100100; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 1974,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110101; i1 = 6'b000101; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110101; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 1975,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011011; i1 = 6'b011010; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011011; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 1976,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011010; i1 = 6'b000010; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011010; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 1977,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001110; i1 = 6'b100001; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001110; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 1978,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100010; i1 = 6'b111010; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100010; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 1979,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111000; i1 = 6'b011010; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111000; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 1980,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011001; i1 = 6'b101111; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011001; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 1981,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b110111; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 1982,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000110; i1 = 6'b010000; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000110; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 1983,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101011; i1 = 6'b101010; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101011; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 1984,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000010; i1 = 6'b111100; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000010; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 1985,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100010; i1 = 6'b110111; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100010; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 1986,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110011; i1 = 6'b111110; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110011; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 1987,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110100; i1 = 6'b000010; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110100; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 1988,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111000; i1 = 6'b111111; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111000; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 1989,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b000010; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 1990,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000000; i1 = 6'b110000; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000000; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 1991,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110110; i1 = 6'b010100; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110110; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 1992,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011100; i1 = 6'b011010; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011100; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 1993,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b001100; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 1994,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000000; i1 = 6'b101001; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000000; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 1995,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111101; i1 = 6'b001010; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111101; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 1996,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b100001; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 1997,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b010101; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 1998,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b000100; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 1999,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111101; i1 = 6'b100101; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111101; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 2000,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101101; i1 = 6'b101001; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101101; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 2001,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001101; i1 = 6'b000011; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001101; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 2002,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010010; i1 = 6'b111011; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010010; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 2003,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101110; i1 = 6'b001101; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101110; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 2004,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b011000; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 2005,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b110011; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 2006,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010000; i1 = 6'b010001; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010000; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 2007,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110110; i1 = 6'b000001; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110110; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 2008,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010101; i1 = 6'b000011; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010101; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 2009,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010000; i1 = 6'b000101; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010000; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 2010,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110110; i1 = 6'b110110; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110110; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 2011,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000010; i1 = 6'b001001; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000010; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 2012,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110001; i1 = 6'b100110; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110001; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 2013,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b000111; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 2014,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110001; i1 = 6'b111001; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110001; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 2015,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b001111; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 2016,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b000001; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 2017,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000010; i1 = 6'b001011; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000010; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 2018,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101110; i1 = 6'b100100; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101110; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 2019,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b000111; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 2020,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100101; i1 = 6'b100011; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100101; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 2021,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b001011; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 2022,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110100; i1 = 6'b010000; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110100; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 2023,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110011; i1 = 6'b010000; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110011; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 2024,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101100; i1 = 6'b000010; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101100; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 2025,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000110; i1 = 6'b011000; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000110; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 2026,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100010; i1 = 6'b101010; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100010; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 2027,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110011; i1 = 6'b110100; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110011; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 2028,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b100010; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 2029,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b111011; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 2030,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000011; i1 = 6'b101101; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000011; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 2031,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100111; i1 = 6'b101100; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100111; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 2032,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010011; i1 = 6'b011111; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010011; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 2033,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000011; i1 = 6'b001110; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000011; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 2034,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b010010; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 2035,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111100; i1 = 6'b101101; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111100; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 2036,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b011110; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 2037,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000010; i1 = 6'b011111; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000010; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 2038,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100111; i1 = 6'b101111; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100111; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 2039,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110000; i1 = 6'b001010; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110000; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 2040,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110101; i1 = 6'b111001; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110101; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 2041,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b011111; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 2042,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b010011; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 2043,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110011; i1 = 6'b100101; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110011; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 2044,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001100; i1 = 6'b110100; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001100; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 2045,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110000; i1 = 6'b001100; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110000; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 2046,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b100010; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 2047,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b101111; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 2048,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001100; i1 = 6'b001000; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001100; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 2049,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b110100; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 2050,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101001; i1 = 6'b101100; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101001; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 2051,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b010010; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 2052,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101000; i1 = 6'b010101; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101000; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 2053,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110011; i1 = 6'b011110; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110011; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 2054,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011001; i1 = 6'b101010; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011001; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 2055,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b100011; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 2056,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b100010; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 2057,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111111; i1 = 6'b000101; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111111; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 2058,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000100; i1 = 6'b100101; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000100; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 2059,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001110; i1 = 6'b000001; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001110; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 2060,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b010001; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 2061,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b100001; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 2062,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110001; i1 = 6'b101100; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110001; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 2063,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001100; i1 = 6'b100110; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001100; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 2064,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101111; i1 = 6'b100101; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101111; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 2065,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011010; i1 = 6'b110011; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011010; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 2066,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b000011; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 2067,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b111110; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 2068,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110101; i1 = 6'b101001; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110101; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 2069,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100111; i1 = 6'b010101; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100111; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 2070,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101000; i1 = 6'b101110; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101000; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 2071,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b011101; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 2072,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111110; i1 = 6'b011101; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111110; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 2073,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b000010; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 2074,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110000; i1 = 6'b110101; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110000; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 2075,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111110; i1 = 6'b111111; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111110; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 2076,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101110; i1 = 6'b100100; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101110; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 2077,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b101101; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 2078,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b100100; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 2079,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b010101; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 2080,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110111; i1 = 6'b110101; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110111; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 2081,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010011; i1 = 6'b011011; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010011; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 2082,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101000; i1 = 6'b110001; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101000; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 2083,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000000; i1 = 6'b100010; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000000; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 2084,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111001; i1 = 6'b100110; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111001; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 2085,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110101; i1 = 6'b001001; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110101; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 2086,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101111; i1 = 6'b000100; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101111; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 2087,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111010; i1 = 6'b011101; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111010; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 2088,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001001; i1 = 6'b111001; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001001; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 2089,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111001; i1 = 6'b000110; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111001; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 2090,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100111; i1 = 6'b010111; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100111; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 2091,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111110; i1 = 6'b000011; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111110; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 2092,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000111; i1 = 6'b011100; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000111; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 2093,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b101000; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 2094,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010100; i1 = 6'b001011; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010100; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 2095,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b001111; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 2096,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b011000; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 2097,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110100; i1 = 6'b100010; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110100; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 2098,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b001011; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 2099,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101100; i1 = 6'b010000; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101100; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 2100,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b101101; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 2101,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b111010; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 2102,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b001100; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 2103,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b100110; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 2104,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001011; i1 = 6'b111000; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001011; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 2105,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110111; i1 = 6'b111010; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110111; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 2106,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110101; i1 = 6'b000000; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110101; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 2107,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110001; i1 = 6'b011010; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110001; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 2108,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011101; i1 = 6'b110011; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011101; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 2109,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010110; i1 = 6'b001011; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010110; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 2110,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101110; i1 = 6'b001100; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101110; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 2111,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b110000; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 2112,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101110; i1 = 6'b111110; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101110; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 2113,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101101; i1 = 6'b000011; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101101; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 2114,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011100; i1 = 6'b101010; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011100; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 2115,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011000; i1 = 6'b110100; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011000; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 2116,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011000; i1 = 6'b010011; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011000; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 2117,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b010010; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 2118,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110011; i1 = 6'b000001; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110011; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 2119,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b000010; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 2120,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001110; i1 = 6'b010010; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001110; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 2121,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b001111; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 2122,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011011; i1 = 6'b101101; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011011; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 2123,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b110100; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 2124,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b010000; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 2125,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110100; i1 = 6'b001101; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110100; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 2126,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111010; i1 = 6'b011001; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111010; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 2127,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110101; i1 = 6'b000010; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110101; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 2128,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100010; i1 = 6'b001100; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100010; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 2129,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110000; i1 = 6'b100101; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110000; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 2130,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b010000; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 2131,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101111; i1 = 6'b011111; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101111; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 2132,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011001; i1 = 6'b000110; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011001; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 2133,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111101; i1 = 6'b001100; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111101; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 2134,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b101111; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 2135,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001111; i1 = 6'b010011; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001111; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 2136,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b010011; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 2137,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b111110; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 2138,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011111; i1 = 6'b010000; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011111; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 2139,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001111; i1 = 6'b111011; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001111; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 2140,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b111011; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 2141,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b100010; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 2142,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b100110; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 2143,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101101; i1 = 6'b110100; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101101; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 2144,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010010; i1 = 6'b010000; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010010; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 2145,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001110; i1 = 6'b001011; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001110; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 2146,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b000011; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 2147,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111010; i1 = 6'b000001; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111010; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 2148,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011110; i1 = 6'b011101; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011110; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 2149,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b001000; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 2150,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001001; i1 = 6'b010100; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001001; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 2151,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101000; i1 = 6'b001101; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101000; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 2152,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111101; i1 = 6'b010000; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111101; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 2153,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b100011; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 2154,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100101; i1 = 6'b011100; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100101; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 2155,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111111; i1 = 6'b011101; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111111; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 2156,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b010010; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 2157,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b110111; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 2158,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101001; i1 = 6'b000010; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101001; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 2159,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110110; i1 = 6'b000000; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110110; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 2160,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b000110; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 2161,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010001; i1 = 6'b011110; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010001; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 2162,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b010100; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 2163,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b011000; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 2164,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111101; i1 = 6'b111111; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111101; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 2165,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101001; i1 = 6'b100011; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101001; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 2166,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000101; i1 = 6'b110100; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000101; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 2167,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011111; i1 = 6'b010100; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011111; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 2168,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b101001; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 2169,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b011100; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 2170,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111010; i1 = 6'b001011; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111010; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 2171,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101000; i1 = 6'b010111; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101000; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 2172,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001110; i1 = 6'b001001; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001110; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 2173,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011010; i1 = 6'b100110; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011010; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 2174,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110111; i1 = 6'b010100; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110111; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 2175,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000111; i1 = 6'b110001; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000111; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 2176,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001111; i1 = 6'b011001; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001111; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 2177,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100100; i1 = 6'b101000; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100100; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 2178,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100110; i1 = 6'b000000; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100110; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 2179,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b010011; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 2180,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000101; i1 = 6'b011100; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000101; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 2181,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b010111; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 2182,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010101; i1 = 6'b011011; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010101; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 2183,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010011; i1 = 6'b111101; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010011; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 2184,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110110; i1 = 6'b111100; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110110; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 2185,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000000; i1 = 6'b001010; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000000; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 2186,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011101; i1 = 6'b010001; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011101; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 2187,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110101; i1 = 6'b001100; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110101; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 2188,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b111100; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 2189,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b011001; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 2190,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b110101; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 2191,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011110; i1 = 6'b101010; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011110; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 2192,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b011001; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 2193,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001000; i1 = 6'b010011; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001000; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 2194,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110100; i1 = 6'b110100; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110100; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 2195,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111110; i1 = 6'b010100; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111110; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 2196,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101111; i1 = 6'b000110; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101111; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 2197,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b011010; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 2198,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011100; i1 = 6'b100101; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011100; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 2199,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111111; i1 = 6'b110100; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111111; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 2200,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111000; i1 = 6'b101100; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111000; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 2201,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b100100; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 2202,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100010; i1 = 6'b010001; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100010; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 2203,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b011111; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 2204,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111001; i1 = 6'b100000; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111001; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 2205,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110001; i1 = 6'b101011; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110001; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 2206,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101101; i1 = 6'b101100; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101101; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 2207,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110001; i1 = 6'b101010; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110001; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 2208,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b100001; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 2209,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110101; i1 = 6'b110000; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110101; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 2210,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b110000; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 2211,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000100; i1 = 6'b001011; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000100; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 2212,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110100; i1 = 6'b100001; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110100; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 2213,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001001; i1 = 6'b001010; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001001; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 2214,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001110; i1 = 6'b101100; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001110; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 2215,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110101; i1 = 6'b001111; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110101; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 2216,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110001; i1 = 6'b111011; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110001; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 2217,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b100000; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 2218,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000011; i1 = 6'b101111; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000011; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 2219,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000100; i1 = 6'b011011; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000100; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 2220,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b111110; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 2221,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110001; i1 = 6'b000010; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110001; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 2222,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011101; i1 = 6'b110101; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011101; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 2223,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b111111; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 2224,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101011; i1 = 6'b010010; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101011; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 2225,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010010; i1 = 6'b000001; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010010; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 2226,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011010; i1 = 6'b000111; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011010; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 2227,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000100; i1 = 6'b000110; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000100; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 2228,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101000; i1 = 6'b111010; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101000; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 2229,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b100001; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 2230,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011010; i1 = 6'b111011; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011010; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 2231,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011011; i1 = 6'b000000; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011011; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 2232,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100100; i1 = 6'b011001; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100100; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 2233,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b000000; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 2234,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100010; i1 = 6'b100011; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100010; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 2235,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011100; i1 = 6'b101110; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011100; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 2236,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110100; i1 = 6'b000100; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110100; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 2237,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001100; i1 = 6'b100000; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001100; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 2238,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101100; i1 = 6'b100000; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101100; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 2239,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001000; i1 = 6'b000101; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001000; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 2240,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001001; i1 = 6'b111010; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001001; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 2241,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b001011; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 2242,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101011; i1 = 6'b000100; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101011; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 2243,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b110000; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 2244,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100100; i1 = 6'b000110; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100100; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 2245,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111101; i1 = 6'b010101; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111101; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 2246,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b110100; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 2247,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b000110; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 2248,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111111; i1 = 6'b110000; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111111; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 2249,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010111; i1 = 6'b000011; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010111; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 2250,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b101110; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 2251,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101011; i1 = 6'b110010; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101011; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 2252,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111111; i1 = 6'b001001; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111111; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 2253,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b110000; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 2254,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110010; i1 = 6'b011101; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110010; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 2255,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011100; i1 = 6'b101101; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011100; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 2256,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100110; i1 = 6'b111110; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100110; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 2257,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010001; i1 = 6'b110001; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010001; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 2258,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101011; i1 = 6'b100000; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101011; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 2259,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b110000; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 2260,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010011; i1 = 6'b100010; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010011; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 2261,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101000; i1 = 6'b101011; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101000; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 2262,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010011; i1 = 6'b101100; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010011; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 2263,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111001; i1 = 6'b011011; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111001; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 2264,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b111011; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 2265,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b000110; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 2266,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b110011; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 2267,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010110; i1 = 6'b011010; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010110; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 2268,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b110111; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 2269,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100111; i1 = 6'b000101; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100111; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 2270,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101101; i1 = 6'b111100; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101101; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 2271,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110000; i1 = 6'b011011; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110000; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 2272,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000100; i1 = 6'b110001; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000100; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 2273,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111111; i1 = 6'b010111; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111111; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 2274,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b010010; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 2275,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010001; i1 = 6'b000000; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010001; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 2276,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110101; i1 = 6'b001011; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110101; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 2277,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111000; i1 = 6'b001110; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111000; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 2278,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000011; i1 = 6'b010000; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000011; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 2279,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011010; i1 = 6'b111111; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011010; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 2280,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b010101; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 2281,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110010; i1 = 6'b110111; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110010; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 2282,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100001; i1 = 6'b111010; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100001; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 2283,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001101; i1 = 6'b001010; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001101; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 2284,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b000000; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 2285,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000011; i1 = 6'b011100; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000011; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 2286,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100100; i1 = 6'b111001; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100100; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 2287,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b001110; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 2288,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011100; i1 = 6'b001000; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011100; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 2289,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111110; i1 = 6'b111011; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111110; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 2290,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b100100; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 2291,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110111; i1 = 6'b100010; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110111; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 2292,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b110000; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 2293,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b100000; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 2294,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110111; i1 = 6'b001101; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110111; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 2295,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001111; i1 = 6'b001100; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001111; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 2296,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b001011; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 2297,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101000; i1 = 6'b001100; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101000; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 2298,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011101; i1 = 6'b100001; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011101; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 2299,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010001; i1 = 6'b011111; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010001; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 2300,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b010101; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 2301,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010111; i1 = 6'b001001; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010111; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 2302,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b010111; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 2303,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111101; i1 = 6'b101100; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111101; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 2304,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011001; i1 = 6'b010101; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011001; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 2305,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b100110; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 2306,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b001011; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 2307,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110101; i1 = 6'b000010; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110101; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 2308,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111110; i1 = 6'b000110; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111110; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 2309,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b101101; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 2310,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100010; i1 = 6'b011101; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100010; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 2311,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110011; i1 = 6'b010011; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110011; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 2312,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111000; i1 = 6'b000001; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111000; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 2313,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111001; i1 = 6'b010111; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111001; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 2314,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000100; i1 = 6'b110110; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000100; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 2315,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001111; i1 = 6'b111000; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001111; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 2316,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b100110; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 2317,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001110; i1 = 6'b111000; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001110; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 2318,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111000; i1 = 6'b101011; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111000; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 2319,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b100000; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 2320,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101001; i1 = 6'b110111; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101001; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 2321,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010100; i1 = 6'b011111; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010100; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 2322,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b100010; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 2323,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010010; i1 = 6'b001010; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010010; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 2324,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001110; i1 = 6'b010110; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001110; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 2325,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100100; i1 = 6'b010010; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100100; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 2326,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010110; i1 = 6'b001100; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010110; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 2327,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b110101; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 2328,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001101; i1 = 6'b111110; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001101; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 2329,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100101; i1 = 6'b000100; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100101; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 2330,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011011; i1 = 6'b100111; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011011; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 2331,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101001; i1 = 6'b111011; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101001; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 2332,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010100; i1 = 6'b110101; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010100; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 2333,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b111111; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 2334,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000101; i1 = 6'b010011; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000101; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 2335,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110100; i1 = 6'b010100; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110100; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 2336,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111010; i1 = 6'b000001; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111010; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 2337,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110100; i1 = 6'b110101; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110100; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 2338,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110011; i1 = 6'b010111; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110011; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 2339,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b001100; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 2340,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101011; i1 = 6'b101001; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101011; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 2341,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000110; i1 = 6'b001000; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000110; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 2342,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000010; i1 = 6'b110000; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000010; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 2343,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001000; i1 = 6'b111001; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001000; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 2344,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b101001; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 2345,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011000; i1 = 6'b101001; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011000; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 2346,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b100001; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 2347,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111110; i1 = 6'b001010; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111110; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 2348,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100001; i1 = 6'b111110; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100001; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 2349,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100001; i1 = 6'b111111; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100001; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 2350,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b011001; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 2351,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111101; i1 = 6'b011111; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111101; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 2352,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011010; i1 = 6'b100101; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011010; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 2353,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110111; i1 = 6'b011000; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110111; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 2354,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100100; i1 = 6'b001000; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100100; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 2355,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b110001; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 2356,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111111; i1 = 6'b110110; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111111; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 2357,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b111010; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 2358,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100010; i1 = 6'b000000; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100010; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 2359,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b110101; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 2360,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100110; i1 = 6'b111010; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100110; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 2361,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000100; i1 = 6'b100110; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000100; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 2362,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101101; i1 = 6'b010110; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101101; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 2363,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b010011; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 2364,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100100; i1 = 6'b100110; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100100; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 2365,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100111; i1 = 6'b101000; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100111; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 2366,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111110; i1 = 6'b001011; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111110; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 2367,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101011; i1 = 6'b111000; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101011; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 2368,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001011; i1 = 6'b011101; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001011; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 2369,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100111; i1 = 6'b100010; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100111; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 2370,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011111; i1 = 6'b011001; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011111; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 2371,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000000; i1 = 6'b011101; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000000; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 2372,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011100; i1 = 6'b100010; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011100; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 2373,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110111; i1 = 6'b000000; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110111; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 2374,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101000; i1 = 6'b000001; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101000; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 2375,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b110100; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 2376,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111101; i1 = 6'b100001; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111101; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 2377,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101001; i1 = 6'b010111; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101001; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 2378,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101011; i1 = 6'b000110; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101011; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 2379,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000111; i1 = 6'b101111; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000111; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 2380,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001110; i1 = 6'b100011; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001110; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 2381,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011100; i1 = 6'b101010; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011100; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 2382,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100110; i1 = 6'b110000; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100110; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 2383,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101001; i1 = 6'b100000; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101001; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 2384,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010001; i1 = 6'b011101; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010001; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 2385,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b101100; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 2386,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b100000; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 2387,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110100; i1 = 6'b010100; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110100; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 2388,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011001; i1 = 6'b010001; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011001; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 2389,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000100; i1 = 6'b000100; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000100; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 2390,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100010; i1 = 6'b111101; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100010; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 2391,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001100; i1 = 6'b101011; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001100; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 2392,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b111100; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 2393,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b110001; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 2394,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101001; i1 = 6'b010001; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101001; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 2395,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000011; i1 = 6'b001011; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000011; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 2396,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101101; i1 = 6'b110111; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101101; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 2397,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010110; i1 = 6'b101100; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010110; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 2398,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b110111; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 2399,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011101; i1 = 6'b110110; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011101; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 2400,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b010110; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 2401,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010001; i1 = 6'b000011; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010001; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 2402,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110011; i1 = 6'b100000; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110011; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 2403,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011010; i1 = 6'b001000; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011010; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 2404,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b111000; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 2405,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b110001; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 2406,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000101; i1 = 6'b110001; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000101; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 2407,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011100; i1 = 6'b100001; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011100; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 2408,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010100; i1 = 6'b101001; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010100; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 2409,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010001; i1 = 6'b010010; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010001; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 2410,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010001; i1 = 6'b101101; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010001; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 2411,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b101101; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 2412,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b010000; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 2413,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101110; i1 = 6'b011100; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101110; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 2414,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000011; i1 = 6'b011111; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000011; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 2415,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100111; i1 = 6'b011111; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100111; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 2416,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011011; i1 = 6'b101110; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011011; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 2417,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010100; i1 = 6'b010101; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010100; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 2418,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101000; i1 = 6'b101101; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101000; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 2419,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010101; i1 = 6'b000011; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010101; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 2420,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001001; i1 = 6'b010101; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001001; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 2421,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100010; i1 = 6'b010000; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100010; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 2422,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100101; i1 = 6'b100101; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100101; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 2423,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001000; i1 = 6'b100101; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001000; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 2424,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010101; i1 = 6'b001001; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010101; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 2425,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000110; i1 = 6'b111110; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000110; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 2426,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110110; i1 = 6'b101101; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110110; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 2427,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b111111; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 2428,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110011; i1 = 6'b010100; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110011; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 2429,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001000; i1 = 6'b101001; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001000; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 2430,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010110; i1 = 6'b101011; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010110; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 2431,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101110; i1 = 6'b111111; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101110; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 2432,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010101; i1 = 6'b000100; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010101; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 2433,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b000100; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 2434,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b101110; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 2435,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b101010; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 2436,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b111010; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 2437,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001001; i1 = 6'b110001; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001001; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 2438,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010100; i1 = 6'b000011; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010100; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 2439,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110011; i1 = 6'b001010; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110011; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 2440,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100100; i1 = 6'b110001; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100100; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 2441,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000101; i1 = 6'b110110; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000101; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 2442,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b110001; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 2443,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011001; i1 = 6'b101110; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011001; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 2444,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001101; i1 = 6'b000000; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001101; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 2445,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b111000; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 2446,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b011100; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 2447,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100011; i1 = 6'b101100; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100011; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 2448,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011011; i1 = 6'b001110; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011011; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 2449,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100001; i1 = 6'b001100; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100001; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 2450,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b001101; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 2451,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b001011; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 2452,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101100; i1 = 6'b010110; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101100; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 2453,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100010; i1 = 6'b001100; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100010; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 2454,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b011100; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 2455,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b010101; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 2456,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010001; i1 = 6'b011000; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010001; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 2457,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011010; i1 = 6'b011001; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011010; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 2458,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000000; i1 = 6'b100111; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000000; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 2459,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001001; i1 = 6'b000010; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001001; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 2460,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101110; i1 = 6'b010101; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101110; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 2461,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101110; i1 = 6'b011011; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101110; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 2462,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b101001; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 2463,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110001; i1 = 6'b101101; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110001; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 2464,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110101; i1 = 6'b011010; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110101; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 2465,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b101100; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 2466,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101011; i1 = 6'b001010; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101011; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 2467,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011111; i1 = 6'b000110; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011111; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 2468,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101110; i1 = 6'b100010; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101110; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 2469,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100101; i1 = 6'b011101; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100101; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 2470,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101101; i1 = 6'b010011; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101101; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 2471,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111000; i1 = 6'b010111; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111000; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 2472,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010110; i1 = 6'b001001; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010110; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 2473,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b000110; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 2474,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111010; i1 = 6'b001100; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111010; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 2475,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111111; i1 = 6'b001011; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111111; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 2476,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b011110; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 2477,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111111; i1 = 6'b001111; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111111; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 2478,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000100; i1 = 6'b000111; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000100; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 2479,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001001; i1 = 6'b001101; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001001; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 2480,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000011; i1 = 6'b100100; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000011; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 2481,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001000; i1 = 6'b000011; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001000; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 2482,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100011; i1 = 6'b000001; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100011; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 2483,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101110; i1 = 6'b010011; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101110; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 2484,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110100; i1 = 6'b000000; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110100; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 2485,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b001000; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 2486,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b000011; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 2487,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b001011; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 2488,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011101; i1 = 6'b001011; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011101; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 2489,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b000011; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 2490,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101011; i1 = 6'b110111; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101011; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 2491,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011011; i1 = 6'b010101; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011011; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 2492,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010001; i1 = 6'b110101; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010001; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 2493,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b111001; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 2494,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001000; i1 = 6'b010001; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001000; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 2495,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100011; i1 = 6'b101001; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100011; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 2496,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010110; i1 = 6'b101110; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010110; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 2497,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b100101; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 2498,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b101101; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 2499,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010110; i1 = 6'b011011; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010110; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 2500,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011010; i1 = 6'b011111; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011010; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 2501,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010110; i1 = 6'b011110; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010110; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 2502,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100101; i1 = 6'b101101; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100101; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 2503,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b001011; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 2504,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b100101; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 2505,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110110; i1 = 6'b101111; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110110; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 2506,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b100110; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 2507,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b010100; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 2508,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000000; i1 = 6'b010110; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000000; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 2509,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b100101; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 2510,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111001; i1 = 6'b101011; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111001; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 2511,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000000; i1 = 6'b110010; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000000; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 2512,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b011011; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 2513,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011101; i1 = 6'b110010; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011101; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 2514,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011011; i1 = 6'b011110; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011011; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 2515,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b011110; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 2516,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b110000; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 2517,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111010; i1 = 6'b110000; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111010; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 2518,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101101; i1 = 6'b101111; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101101; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 2519,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111000; i1 = 6'b000101; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111000; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 2520,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b110000; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 2521,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110110; i1 = 6'b010000; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110110; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 2522,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b100010; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 2523,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110000; i1 = 6'b110110; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110000; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 2524,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010110; i1 = 6'b000011; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010110; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 2525,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010001; i1 = 6'b111011; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010001; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 2526,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100001; i1 = 6'b001011; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100001; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 2527,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b000000; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 2528,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b001101; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 2529,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110001; i1 = 6'b011100; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110001; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 2530,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b011110; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 2531,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010110; i1 = 6'b111010; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010110; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 2532,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110010; i1 = 6'b101011; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110010; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 2533,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111110; i1 = 6'b101001; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111110; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 2534,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110011; i1 = 6'b101010; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110011; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 2535,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b001010; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 2536,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b100110; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 2537,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b111110; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 2538,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b111110; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 2539,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110001; i1 = 6'b100001; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110001; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 2540,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111001; i1 = 6'b111111; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111001; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 2541,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011100; i1 = 6'b100100; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011100; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 2542,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000010; i1 = 6'b100100; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000010; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 2543,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111111; i1 = 6'b101101; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111111; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 2544,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010101; i1 = 6'b001011; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010101; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 2545,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101011; i1 = 6'b001110; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101011; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 2546,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000000; i1 = 6'b111101; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000000; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 2547,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b101010; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 2548,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111110; i1 = 6'b110011; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111110; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 2549,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b111101; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 2550,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000100; i1 = 6'b001001; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000100; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 2551,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b011100; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 2552,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b000111; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 2553,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100111; i1 = 6'b010001; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100111; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 2554,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001110; i1 = 6'b101000; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001110; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 2555,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100001; i1 = 6'b010000; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100001; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 2556,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000111; i1 = 6'b101110; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000111; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 2557,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b110110; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 2558,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100001; i1 = 6'b001000; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100001; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 2559,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b000111; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 2560,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010001; i1 = 6'b010111; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010001; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 2561,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b100011; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 2562,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011011; i1 = 6'b110101; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011011; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 2563,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111010; i1 = 6'b110111; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111010; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 2564,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b000111; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 2565,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110010; i1 = 6'b101001; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110010; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 2566,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110010; i1 = 6'b101100; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110010; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 2567,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111101; i1 = 6'b011010; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111101; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 2568,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010111; i1 = 6'b110101; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010111; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 2569,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101000; i1 = 6'b001110; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101000; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 2570,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b011001; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 2571,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100010; i1 = 6'b010010; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100010; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 2572,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111010; i1 = 6'b011011; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111010; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 2573,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111110; i1 = 6'b101010; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111110; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 2574,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b100101; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 2575,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b110000; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 2576,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101100; i1 = 6'b011100; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101100; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 2577,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110001; i1 = 6'b100100; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110001; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 2578,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101111; i1 = 6'b111101; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101111; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 2579,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101001; i1 = 6'b001101; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101001; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 2580,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000111; i1 = 6'b101011; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000111; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 2581,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000101; i1 = 6'b111010; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000101; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 2582,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001000; i1 = 6'b111010; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001000; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 2583,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100111; i1 = 6'b110000; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100111; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 2584,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011011; i1 = 6'b000101; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011011; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 2585,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111101; i1 = 6'b111111; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111101; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 2586,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000101; i1 = 6'b010111; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000101; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 2587,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011001; i1 = 6'b100000; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011001; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 2588,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001001; i1 = 6'b010111; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001001; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 2589,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011011; i1 = 6'b111010; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011011; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 2590,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111000; i1 = 6'b000100; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111000; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 2591,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001100; i1 = 6'b010010; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001100; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 2592,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b001101; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 2593,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000100; i1 = 6'b100010; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000100; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 2594,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110111; i1 = 6'b000001; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110111; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 2595,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110101; i1 = 6'b000110; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110101; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 2596,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101001; i1 = 6'b100011; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101001; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 2597,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111110; i1 = 6'b010011; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111110; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 2598,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b100011; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 2599,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011110; i1 = 6'b000010; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011110; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 2600,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b010000; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 2601,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010011; i1 = 6'b000101; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010011; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 2602,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110111; i1 = 6'b011110; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110111; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 2603,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b011011; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 2604,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b000010; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 2605,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011010; i1 = 6'b010100; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011010; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 2606,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100010; i1 = 6'b110110; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100010; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 2607,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b100001; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 2608,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110101; i1 = 6'b101010; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110101; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 2609,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b100100; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 2610,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101110; i1 = 6'b111111; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101110; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 2611,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111010; i1 = 6'b111010; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111010; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 2612,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011011; i1 = 6'b011101; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011011; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 2613,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111000; i1 = 6'b010111; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111000; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 2614,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000000; i1 = 6'b110110; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000000; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 2615,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100100; i1 = 6'b100001; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100100; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 2616,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111111; i1 = 6'b111110; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111111; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 2617,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111101; i1 = 6'b000100; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111101; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 2618,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101110; i1 = 6'b010101; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101110; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 2619,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101100; i1 = 6'b010100; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101100; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 2620,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110011; i1 = 6'b110000; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110011; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 2621,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010111; i1 = 6'b100110; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010111; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 2622,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001001; i1 = 6'b011101; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001001; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 2623,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101001; i1 = 6'b000110; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101001; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 2624,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110110; i1 = 6'b110011; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110110; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 2625,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b011100; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 2626,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011010; i1 = 6'b000101; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011010; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 2627,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001100; i1 = 6'b010000; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001100; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 2628,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010111; i1 = 6'b110000; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010111; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 2629,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011000; i1 = 6'b111000; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011000; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 2630,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010000; i1 = 6'b010000; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010000; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 2631,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b100010; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 2632,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b011111; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 2633,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011011; i1 = 6'b100010; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011011; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 2634,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b110000; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 2635,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110111; i1 = 6'b000011; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110111; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 2636,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101011; i1 = 6'b011000; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101011; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 2637,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010001; i1 = 6'b100111; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010001; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 2638,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001101; i1 = 6'b110000; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001101; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 2639,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011110; i1 = 6'b010010; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011110; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 2640,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b100100; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 2641,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000110; i1 = 6'b111011; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000110; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 2642,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000011; i1 = 6'b011101; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000011; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 2643,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111111; i1 = 6'b001010; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111111; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 2644,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b001110; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 2645,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001011; i1 = 6'b100110; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001011; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 2646,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110011; i1 = 6'b110001; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110011; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 2647,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000111; i1 = 6'b101110; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000111; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 2648,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000110; i1 = 6'b011010; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000110; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 2649,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b100001; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 2650,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011011; i1 = 6'b000100; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011011; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 2651,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010001; i1 = 6'b001111; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010001; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 2652,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b110001; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 2653,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100010; i1 = 6'b000111; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100010; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 2654,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000011; i1 = 6'b000001; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000011; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 2655,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000110; i1 = 6'b101101; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000110; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 2656,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001110; i1 = 6'b000110; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001110; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 2657,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001110; i1 = 6'b000001; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001110; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 2658,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b001100; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 2659,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011001; i1 = 6'b101100; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011001; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 2660,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010001; i1 = 6'b100010; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010001; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 2661,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101001; i1 = 6'b011111; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101001; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 2662,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011110; i1 = 6'b110110; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011110; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 2663,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b101010; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 2664,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101000; i1 = 6'b101001; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101000; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 2665,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110000; i1 = 6'b111111; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110000; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 2666,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000100; i1 = 6'b111111; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000100; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 2667,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000100; i1 = 6'b011100; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000100; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 2668,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111010; i1 = 6'b111101; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111010; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 2669,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000000; i1 = 6'b000100; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000000; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 2670,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000000; i1 = 6'b000010; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000000; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 2671,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101101; i1 = 6'b000010; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101101; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 2672,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b010101; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 2673,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001000; i1 = 6'b100110; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001000; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 2674,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111110; i1 = 6'b000111; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111110; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 2675,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111110; i1 = 6'b101000; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111110; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 2676,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011010; i1 = 6'b011100; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011010; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 2677,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010110; i1 = 6'b111101; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010110; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 2678,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010100; i1 = 6'b111011; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010100; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 2679,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000000; i1 = 6'b010010; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000000; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 2680,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111000; i1 = 6'b010001; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111000; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 2681,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001101; i1 = 6'b110111; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001101; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 2682,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b000010; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 2683,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010101; i1 = 6'b111101; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010101; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 2684,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b100001; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 2685,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111110; i1 = 6'b111110; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111110; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 2686,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111000; i1 = 6'b110111; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111000; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 2687,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011101; i1 = 6'b111110; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011101; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 2688,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000100; i1 = 6'b110010; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000100; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 2689,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010001; i1 = 6'b111010; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010001; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 2690,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110101; i1 = 6'b101111; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110101; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 2691,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b101101; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 2692,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b001101; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 2693,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001011; i1 = 6'b010010; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001011; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 2694,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011001; i1 = 6'b110010; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011001; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 2695,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011101; i1 = 6'b101101; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011101; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 2696,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b010011; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 2697,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001000; i1 = 6'b110100; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001000; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 2698,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b111101; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 2699,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101001; i1 = 6'b000100; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101001; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 2700,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011010; i1 = 6'b101001; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011010; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 2701,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011100; i1 = 6'b011111; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011100; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 2702,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b111010; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 2703,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101100; i1 = 6'b001110; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101100; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 2704,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011011; i1 = 6'b000100; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011011; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 2705,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101101; i1 = 6'b011111; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101101; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 2706,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b111001; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 2707,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010101; i1 = 6'b110010; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010101; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 2708,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010101; i1 = 6'b110001; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010101; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 2709,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100111; i1 = 6'b001111; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100111; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 2710,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b011000; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 2711,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011101; i1 = 6'b110001; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011101; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 2712,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000100; i1 = 6'b000010; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000100; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 2713,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b001001; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 2714,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b010111; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 2715,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b100000; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 2716,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010100; i1 = 6'b100010; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010100; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 2717,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100101; i1 = 6'b100111; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100101; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 2718,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000111; i1 = 6'b011111; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000111; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 2719,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b001010; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 2720,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b010011; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 2721,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011010; i1 = 6'b100100; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011010; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 2722,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010110; i1 = 6'b101000; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010110; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 2723,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000110; i1 = 6'b010001; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000110; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 2724,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010100; i1 = 6'b111100; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010100; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 2725,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110110; i1 = 6'b111010; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110110; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 2726,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010111; i1 = 6'b001000; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010111; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 2727,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b110000; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 2728,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010001; i1 = 6'b100100; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010001; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 2729,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b110010; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 2730,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110010; i1 = 6'b001111; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110010; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 2731,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101111; i1 = 6'b111010; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101111; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 2732,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010001; i1 = 6'b001111; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010001; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 2733,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000110; i1 = 6'b000011; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000110; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 2734,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000000; i1 = 6'b001001; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000000; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 2735,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010110; i1 = 6'b010010; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010110; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 2736,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100101; i1 = 6'b100010; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100101; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 2737,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011001; i1 = 6'b000111; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011001; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 2738,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000011; i1 = 6'b010100; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000011; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 2739,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000101; i1 = 6'b100000; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000101; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 2740,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000101; i1 = 6'b111111; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000101; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 2741,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b000111; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 2742,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010100; i1 = 6'b110001; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010100; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 2743,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110000; i1 = 6'b011001; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110000; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 2744,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110100; i1 = 6'b011101; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110100; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 2745,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011001; i1 = 6'b001110; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011001; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 2746,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001001; i1 = 6'b001110; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001001; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 2747,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b000010; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 2748,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010101; i1 = 6'b111111; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010101; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 2749,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100101; i1 = 6'b000110; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100101; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 2750,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b010100; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 2751,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110001; i1 = 6'b011111; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110001; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 2752,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100001; i1 = 6'b100000; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100001; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 2753,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001100; i1 = 6'b011110; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001100; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 2754,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101100; i1 = 6'b100111; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101100; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 2755,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001001; i1 = 6'b110111; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001001; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 2756,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110110; i1 = 6'b000110; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110110; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 2757,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b111101; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 2758,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b111000; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 2759,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010111; i1 = 6'b010111; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010111; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 2760,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111101; i1 = 6'b100010; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111101; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 2761,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b001101; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 2762,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001011; i1 = 6'b111101; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001011; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 2763,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100001; i1 = 6'b010011; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100001; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 2764,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011111; i1 = 6'b010011; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011111; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 2765,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b100111; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 2766,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100010; i1 = 6'b011001; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100010; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 2767,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100100; i1 = 6'b101001; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100100; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 2768,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b101011; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 2769,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b111100; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 2770,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b100100; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 2771,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111101; i1 = 6'b010001; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111101; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 2772,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100001; i1 = 6'b101001; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100001; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 2773,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001101; i1 = 6'b101011; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001101; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 2774,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011100; i1 = 6'b011100; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011100; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 2775,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011001; i1 = 6'b100101; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011001; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 2776,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010001; i1 = 6'b100101; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010001; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 2777,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011000; i1 = 6'b000000; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011000; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 2778,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101111; i1 = 6'b100010; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101111; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 2779,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010101; i1 = 6'b111100; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010101; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 2780,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110100; i1 = 6'b001111; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110100; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 2781,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110100; i1 = 6'b000001; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110100; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 2782,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000011; i1 = 6'b010111; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000011; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 2783,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000101; i1 = 6'b001111; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000101; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 2784,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101011; i1 = 6'b001000; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101011; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 2785,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b111110; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 2786,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110100; i1 = 6'b110100; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110100; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 2787,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010111; i1 = 6'b110010; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010111; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 2788,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111001; i1 = 6'b111100; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111001; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 2789,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100000; i1 = 6'b001011; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100000; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 2790,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b001110; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 2791,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b000111; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 2792,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b011011; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 2793,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b001101; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 2794,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110001; i1 = 6'b110001; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110001; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 2795,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001110; i1 = 6'b100010; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001110; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 2796,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110001; i1 = 6'b010011; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110001; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 2797,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b101101; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 2798,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000000; i1 = 6'b001100; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000000; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 2799,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b110110; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 2800,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011101; i1 = 6'b100000; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011101; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 2801,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b110111; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 2802,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010101; i1 = 6'b001100; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010101; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 2803,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100111; i1 = 6'b010011; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100111; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 2804,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111110; i1 = 6'b011011; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111110; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 2805,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b011011; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 2806,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b101001; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 2807,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b101011; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 2808,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010101; i1 = 6'b010011; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010101; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 2809,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b010011; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 2810,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010101; i1 = 6'b100011; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010101; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 2811,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100100; i1 = 6'b110000; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100100; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 2812,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001110; i1 = 6'b110001; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001110; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 2813,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111111; i1 = 6'b101101; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111111; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 2814,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000110; i1 = 6'b101100; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000110; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 2815,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b001100; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 2816,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011110; i1 = 6'b110000; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011110; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 2817,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000100; i1 = 6'b001010; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000100; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 2818,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011001; i1 = 6'b010000; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011001; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 2819,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100001; i1 = 6'b001010; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100001; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 2820,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011010; i1 = 6'b110010; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011010; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 2821,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110000; i1 = 6'b011110; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110000; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 2822,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101011; i1 = 6'b111111; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101011; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 2823,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110011; i1 = 6'b011000; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110011; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 2824,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b101110; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 2825,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b011010; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 2826,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011011; i1 = 6'b010111; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011011; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 2827,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b101001; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 2828,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110101; i1 = 6'b001101; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110101; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 2829,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b000100; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 2830,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101110; i1 = 6'b101001; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101110; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 2831,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b011101; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 2832,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b011001; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 2833,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011010; i1 = 6'b001101; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011010; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 2834,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100000; i1 = 6'b001000; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100000; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 2835,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001110; i1 = 6'b110110; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001110; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 2836,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b100000; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 2837,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b110001; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 2838,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011011; i1 = 6'b001111; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011011; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 2839,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b111110; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 2840,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b110111; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 2841,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110100; i1 = 6'b101111; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110100; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 2842,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001100; i1 = 6'b100100; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001100; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 2843,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001000; i1 = 6'b101000; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001000; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 2844,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110100; i1 = 6'b000101; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110100; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 2845,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110000; i1 = 6'b000101; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110000; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 2846,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111010; i1 = 6'b111100; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111010; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 2847,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b010110; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 2848,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111101; i1 = 6'b011001; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111101; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 2849,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101110; i1 = 6'b011111; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101110; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 2850,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101101; i1 = 6'b101110; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101101; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 2851,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001110; i1 = 6'b111100; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001110; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 2852,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101110; i1 = 6'b010001; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101110; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 2853,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111010; i1 = 6'b101100; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111010; i1 = 6'b101100; | Outputs: sum=%b | Expected: sum=%d",
                 2854,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110101; i1 = 6'b011001; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110101; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 2855,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000011; i1 = 6'b110010; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000011; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 2856,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110111; i1 = 6'b001100; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110111; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 2857,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010110; i1 = 6'b101101; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010110; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 2858,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b001111; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 2859,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100010; i1 = 6'b100100; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100010; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 2860,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100110; i1 = 6'b000010; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100110; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 2861,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101101; i1 = 6'b110010; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101101; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 2862,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100010; i1 = 6'b010101; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100010; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 2863,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011101; i1 = 6'b110001; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011101; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 2864,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b101000; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 2865,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100010; i1 = 6'b101001; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100010; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 2866,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111000; i1 = 6'b011011; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111000; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 2867,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000010; i1 = 6'b000011; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000010; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 2868,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b010001; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 2869,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b101111; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 2870,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101000; i1 = 6'b011011; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101000; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 2871,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100001; i1 = 6'b101101; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100001; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 2872,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010111; i1 = 6'b000001; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010111; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 2873,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000101; i1 = 6'b011101; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000101; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 2874,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110000; i1 = 6'b001011; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110000; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 2875,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b110110; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 2876,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011100; i1 = 6'b010101; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011100; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 2877,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b110100; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 2878,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101100; i1 = 6'b011011; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101100; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 2879,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110011; i1 = 6'b000000; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110011; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 2880,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b000101; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 2881,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001011; i1 = 6'b101101; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001011; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 2882,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100010; i1 = 6'b101110; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100010; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 2883,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b000011; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 2884,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100010; i1 = 6'b001111; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100010; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 2885,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111110; i1 = 6'b100111; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111110; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 2886,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000000; i1 = 6'b011100; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000000; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 2887,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010010; i1 = 6'b111010; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010010; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 2888,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b111100; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 2889,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110110; i1 = 6'b101001; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110110; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 2890,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011010; i1 = 6'b010000; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011010; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 2891,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010011; i1 = 6'b100100; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010011; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 2892,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b011110; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b011110; | Outputs: sum=%b | Expected: sum=%d",
                 2893,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000111; i1 = 6'b110011; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000111; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 2894,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b001011; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 2895,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000000; i1 = 6'b101111; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000000; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 2896,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111000; i1 = 6'b100001; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111000; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 2897,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100010; i1 = 6'b011111; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100010; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 2898,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111110; i1 = 6'b110111; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111110; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 2899,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b100111; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 2900,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110011; i1 = 6'b110010; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110011; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 2901,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b111101; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 2902,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000111; i1 = 6'b000101; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000111; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 2903,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b000111; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 2904,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101101; i1 = 6'b100100; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101101; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 2905,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110011; i1 = 6'b010010; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110011; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 2906,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010000; i1 = 6'b110110; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010000; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 2907,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000111; i1 = 6'b001000; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000111; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 2908,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111111; i1 = 6'b100001; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111111; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 2909,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011100; i1 = 6'b111100; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011100; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 2910,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000110; i1 = 6'b100110; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000110; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 2911,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010001; i1 = 6'b001001; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010001; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 2912,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011010; i1 = 6'b100110; // Expected: {'sum': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011010; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 2913,
                 
                 sum
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111101; i1 = 6'b001000; // Expected: {'sum': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111101; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 2914,
                 
                 sum
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b100010; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 2915,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011011; i1 = 6'b101000; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011011; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 2916,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110011; i1 = 6'b011010; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110011; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 2917,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b110101; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 2918,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110101; i1 = 6'b011011; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110101; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 2919,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000111; i1 = 6'b011010; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000111; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 2920,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000110; i1 = 6'b100111; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000110; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 2921,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010011; i1 = 6'b010100; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010011; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 2922,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010111; i1 = 6'b001010; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010111; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 2923,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000100; i1 = 6'b101110; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000100; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 2924,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b101111; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 2925,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b000011; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 2926,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100001; i1 = 6'b010101; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100001; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 2927,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b111110; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 2928,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b011011; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 2929,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101011; i1 = 6'b111101; // Expected: {'sum': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101011; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 2930,
                 
                 sum
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110010; i1 = 6'b011011; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110010; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 2931,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101000; i1 = 6'b101001; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101000; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 2932,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010101; i1 = 6'b100100; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010101; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 2933,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110111; i1 = 6'b111100; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110111; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 2934,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b111010; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 2935,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011100; i1 = 6'b101000; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011100; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 2936,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b000110; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 2937,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010010; i1 = 6'b010001; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010010; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 2938,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100001; i1 = 6'b000110; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100001; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 2939,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011000; i1 = 6'b011001; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011000; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 2940,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b110000; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 2941,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001000; i1 = 6'b101010; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001000; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 2942,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010011; i1 = 6'b110001; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010011; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 2943,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001001; i1 = 6'b001001; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001001; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 2944,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110011; i1 = 6'b110011; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110011; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 2945,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111111; i1 = 6'b011010; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111111; i1 = 6'b011010; | Outputs: sum=%b | Expected: sum=%d",
                 2946,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000110; i1 = 6'b001100; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000110; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 2947,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011011; i1 = 6'b001101; // Expected: {'sum': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011011; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 2948,
                 
                 sum
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110001; i1 = 6'b101001; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110001; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 2949,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010000; i1 = 6'b011011; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010000; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 2950,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b111001; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 2951,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110110; i1 = 6'b001100; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110110; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 2952,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100100; i1 = 6'b100000; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100100; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 2953,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000110; i1 = 6'b101011; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000110; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 2954,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001111; i1 = 6'b010101; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001111; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 2955,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100100; i1 = 6'b110101; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100100; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 2956,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111111; i1 = 6'b100010; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111111; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 2957,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111111; i1 = 6'b100111; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111111; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 2958,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101011; i1 = 6'b101000; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101011; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 2959,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b011001; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 2960,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110000; i1 = 6'b110110; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110000; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 2961,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100100; i1 = 6'b000110; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100100; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 2962,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b010110; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 2963,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111111; i1 = 6'b011000; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111111; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 2964,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100101; i1 = 6'b101000; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100101; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 2965,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101001; i1 = 6'b101000; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101001; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 2966,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000010; i1 = 6'b110011; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000010; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 2967,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001011; i1 = 6'b000011; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001011; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 2968,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b100010; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 2969,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011010; i1 = 6'b010010; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011010; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 2970,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011101; i1 = 6'b001001; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011101; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 2971,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111001; i1 = 6'b100101; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111001; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 2972,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000011; i1 = 6'b001100; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000011; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 2973,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100001; i1 = 6'b000111; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100001; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 2974,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000100; i1 = 6'b001000; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000100; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 2975,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000100; i1 = 6'b111011; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000100; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 2976,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000010; i1 = 6'b011011; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000010; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 2977,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111101; i1 = 6'b110001; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111101; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 2978,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b111111; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 2979,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010000; i1 = 6'b000000; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010000; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 2980,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100001; i1 = 6'b100001; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100001; i1 = 6'b100001; | Outputs: sum=%b | Expected: sum=%d",
                 2981,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011011; i1 = 6'b010010; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011011; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 2982,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b001010; // Expected: {'sum': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 2983,
                 
                 sum
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001000; i1 = 6'b111000; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001000; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 2984,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011100; i1 = 6'b110001; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011100; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 2985,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110111; i1 = 6'b001011; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110111; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 2986,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010010; i1 = 6'b111111; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010010; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 2987,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011100; i1 = 6'b110110; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011100; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 2988,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011101; i1 = 6'b000010; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011101; i1 = 6'b000010; | Outputs: sum=%b | Expected: sum=%d",
                 2989,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111010; i1 = 6'b111000; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111010; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 2990,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111100; i1 = 6'b110011; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111100; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 2991,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110101; i1 = 6'b110001; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110101; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 2992,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110100; i1 = 6'b111000; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110100; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 2993,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101100; i1 = 6'b011001; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101100; i1 = 6'b011001; | Outputs: sum=%b | Expected: sum=%d",
                 2994,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b100011; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 2995,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b000001; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b000001; | Outputs: sum=%b | Expected: sum=%d",
                 2996,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000011; i1 = 6'b110100; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000011; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 2997,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001110; i1 = 6'b101001; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001110; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 2998,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000111; i1 = 6'b001110; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000111; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 2999,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111010; i1 = 6'b001000; // Expected: {'sum': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111010; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 3000,
                 
                 sum
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b111101; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b111101; | Outputs: sum=%b | Expected: sum=%d",
                 3001,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000111; i1 = 6'b110010; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000111; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 3002,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110101; i1 = 6'b010000; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110101; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 3003,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110010; i1 = 6'b100110; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110010; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 3004,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111101; i1 = 6'b101001; // Expected: {'sum': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111101; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 3005,
                 
                 sum
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111000; i1 = 6'b000000; // Expected: {'sum': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111000; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 3006,
                 
                 sum
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b010110; // Expected: {'sum': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 3007,
                 
                 sum
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000000; i1 = 6'b001001; // Expected: {'sum': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000000; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 3008,
                 
                 sum
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000110; i1 = 6'b010011; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000110; i1 = 6'b010011; | Outputs: sum=%b | Expected: sum=%d",
                 3009,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000101; i1 = 6'b010010; // Expected: {'sum': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000101; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 3010,
                 
                 sum
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011000; i1 = 6'b010111; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011000; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 3011,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b110010; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 3012,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110111; i1 = 6'b110001; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110111; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 3013,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101000; i1 = 6'b001001; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101000; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 3014,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110010; i1 = 6'b111111; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110010; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 3015,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011010; i1 = 6'b110111; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011010; i1 = 6'b110111; | Outputs: sum=%b | Expected: sum=%d",
                 3016,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101011; i1 = 6'b010001; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101011; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 3017,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001111; i1 = 6'b011100; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001111; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 3018,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111110; i1 = 6'b100011; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111110; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 3019,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001000; i1 = 6'b010010; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001000; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 3020,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b101011; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 3021,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b000110; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 3022,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010111; i1 = 6'b010010; // Expected: {'sum': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010111; i1 = 6'b010010; | Outputs: sum=%b | Expected: sum=%d",
                 3023,
                 
                 sum
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111000; i1 = 6'b101110; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111000; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 3024,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001110; i1 = 6'b010001; // Expected: {'sum': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001110; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 3025,
                 
                 sum
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111011; i1 = 6'b101111; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111011; i1 = 6'b101111; | Outputs: sum=%b | Expected: sum=%d",
                 3026,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000100; i1 = 6'b011111; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000100; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 3027,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b110000; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 3028,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011101; i1 = 6'b110101; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011101; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 3029,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b001000; // Expected: {'sum': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b001000; | Outputs: sum=%b | Expected: sum=%d",
                 3030,
                 
                 sum
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100101; i1 = 6'b111110; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100101; i1 = 6'b111110; | Outputs: sum=%b | Expected: sum=%d",
                 3031,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011111; i1 = 6'b100111; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011111; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 3032,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110011; i1 = 6'b010100; // Expected: {'sum': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110011; i1 = 6'b010100; | Outputs: sum=%b | Expected: sum=%d",
                 3033,
                 
                 sum
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b010101; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 3034,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101110; i1 = 6'b001110; // Expected: {'sum': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101110; i1 = 6'b001110; | Outputs: sum=%b | Expected: sum=%d",
                 3035,
                 
                 sum
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010110; i1 = 6'b100111; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010110; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 3036,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101010; i1 = 6'b010101; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101010; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 3037,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100110; i1 = 6'b111001; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100110; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 3038,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010110; i1 = 6'b100100; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010110; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 3039,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001100; i1 = 6'b111001; // Expected: {'sum': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001100; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 3040,
                 
                 sum
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100111; i1 = 6'b111001; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100111; i1 = 6'b111001; | Outputs: sum=%b | Expected: sum=%d",
                 3041,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101011; i1 = 6'b000000; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101011; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 3042,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111101; i1 = 6'b000101; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111101; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 3043,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111011; i1 = 6'b110001; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111011; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 3044,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010001; i1 = 6'b111011; // Expected: {'sum': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010001; i1 = 6'b111011; | Outputs: sum=%b | Expected: sum=%d",
                 3045,
                 
                 sum
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100110; i1 = 6'b111111; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100110; i1 = 6'b111111; | Outputs: sum=%b | Expected: sum=%d",
                 3046,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010100; i1 = 6'b110101; // Expected: {'sum': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010100; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 3047,
                 
                 sum
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101010; i1 = 6'b000111; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101010; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 3048,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111110; i1 = 6'b111010; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111110; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 3049,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011100; i1 = 6'b110101; // Expected: {'sum': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011100; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 3050,
                 
                 sum
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000001; i1 = 6'b110110; // Expected: {'sum': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000001; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 3051,
                 
                 sum
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100010; i1 = 6'b010101; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100010; i1 = 6'b010101; | Outputs: sum=%b | Expected: sum=%d",
                 3052,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101110; i1 = 6'b010001; // Expected: {'sum': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101110; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 3053,
                 
                 sum
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101000; i1 = 6'b010001; // Expected: {'sum': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101000; i1 = 6'b010001; | Outputs: sum=%b | Expected: sum=%d",
                 3054,
                 
                 sum
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b000000; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b000000; | Outputs: sum=%b | Expected: sum=%d",
                 3055,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000011; i1 = 6'b011000; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000011; i1 = 6'b011000; | Outputs: sum=%b | Expected: sum=%d",
                 3056,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101101; i1 = 6'b111100; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101101; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 3057,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100100; i1 = 6'b100010; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100100; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 3058,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b000001; i1 = 6'b010111; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b000001; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 3059,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100001; i1 = 6'b111100; // Expected: {'sum': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100001; i1 = 6'b111100; | Outputs: sum=%b | Expected: sum=%d",
                 3060,
                 
                 sum
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001100; i1 = 6'b111010; // Expected: {'sum': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001100; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 3061,
                 
                 sum
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001101; i1 = 6'b100100; // Expected: {'sum': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001101; i1 = 6'b100100; | Outputs: sum=%b | Expected: sum=%d",
                 3062,
                 
                 sum
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001110; i1 = 6'b100111; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001110; i1 = 6'b100111; | Outputs: sum=%b | Expected: sum=%d",
                 3063,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b001001; // Expected: {'sum': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 3064,
                 
                 sum
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b001111; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 3065,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011101; i1 = 6'b101000; // Expected: {'sum': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011101; i1 = 6'b101000; | Outputs: sum=%b | Expected: sum=%d",
                 3066,
                 
                 sum
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111111; i1 = 6'b000101; // Expected: {'sum': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111111; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 3067,
                 
                 sum
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001001; i1 = 6'b001111; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001001; i1 = 6'b001111; | Outputs: sum=%b | Expected: sum=%d",
                 3068,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011011; i1 = 6'b110010; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011011; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 3069,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001011; i1 = 6'b001010; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001011; i1 = 6'b001010; | Outputs: sum=%b | Expected: sum=%d",
                 3070,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111111; i1 = 6'b110000; // Expected: {'sum': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111111; i1 = 6'b110000; | Outputs: sum=%b | Expected: sum=%d",
                 3071,
                 
                 sum
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110000; i1 = 6'b110001; // Expected: {'sum': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110000; i1 = 6'b110001; | Outputs: sum=%b | Expected: sum=%d",
                 3072,
                 
                 sum
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000010; i1 = 6'b100110; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000010; i1 = 6'b100110; | Outputs: sum=%b | Expected: sum=%d",
                 3073,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001110; i1 = 6'b111010; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001110; i1 = 6'b111010; | Outputs: sum=%b | Expected: sum=%d",
                 3074,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111110; i1 = 6'b101110; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111110; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 3075,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111100; i1 = 6'b110010; // Expected: {'sum': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111100; i1 = 6'b110010; | Outputs: sum=%b | Expected: sum=%d",
                 3076,
                 
                 sum
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010010; i1 = 6'b000011; // Expected: {'sum': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010010; i1 = 6'b000011; | Outputs: sum=%b | Expected: sum=%d",
                 3077,
                 
                 sum
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111100; i1 = 6'b100000; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111100; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 3078,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001010; i1 = 6'b001011; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001010; i1 = 6'b001011; | Outputs: sum=%b | Expected: sum=%d",
                 3079,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001010; i1 = 6'b100000; // Expected: {'sum': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001010; i1 = 6'b100000; | Outputs: sum=%b | Expected: sum=%d",
                 3080,
                 
                 sum
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101110; i1 = 6'b010110; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101110; i1 = 6'b010110; | Outputs: sum=%b | Expected: sum=%d",
                 3081,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100111; i1 = 6'b110100; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100111; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 3082,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b000110; i1 = 6'b011100; // Expected: {'sum': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b000110; i1 = 6'b011100; | Outputs: sum=%b | Expected: sum=%d",
                 3083,
                 
                 sum
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010110; i1 = 6'b110101; // Expected: {'sum': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010110; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 3084,
                 
                 sum
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001000; i1 = 6'b101110; // Expected: {'sum': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001000; i1 = 6'b101110; | Outputs: sum=%b | Expected: sum=%d",
                 3085,
                 
                 sum
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110111; i1 = 6'b000100; // Expected: {'sum': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110111; i1 = 6'b000100; | Outputs: sum=%b | Expected: sum=%d",
                 3086,
                 
                 sum
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100001; i1 = 6'b011101; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100001; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 3087,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101111; i1 = 6'b100010; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101111; i1 = 6'b100010; | Outputs: sum=%b | Expected: sum=%d",
                 3088,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001100; i1 = 6'b000110; // Expected: {'sum': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001100; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 3089,
                 
                 sum
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001110; i1 = 6'b110011; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001110; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 3090,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101100; i1 = 6'b101001; // Expected: {'sum': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101100; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 3091,
                 
                 sum
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010000; i1 = 6'b100011; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010000; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 3092,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110101; i1 = 6'b101011; // Expected: {'sum': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110101; i1 = 6'b101011; | Outputs: sum=%b | Expected: sum=%d",
                 3093,
                 
                 sum
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011001; i1 = 6'b110110; // Expected: {'sum': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011001; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 3094,
                 
                 sum
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101110; i1 = 6'b010000; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101110; i1 = 6'b010000; | Outputs: sum=%b | Expected: sum=%d",
                 3095,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010101; i1 = 6'b101001; // Expected: {'sum': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010101; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 3096,
                 
                 sum
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b111110; i1 = 6'b010111; // Expected: {'sum': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b111110; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 3097,
                 
                 sum
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110110; i1 = 6'b111000; // Expected: {'sum': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110110; i1 = 6'b111000; | Outputs: sum=%b | Expected: sum=%d",
                 3098,
                 
                 sum
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001110; i1 = 6'b011101; // Expected: {'sum': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001110; i1 = 6'b011101; | Outputs: sum=%b | Expected: sum=%d",
                 3099,
                 
                 sum
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110001; i1 = 6'b110011; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110001; i1 = 6'b110011; | Outputs: sum=%b | Expected: sum=%d",
                 3100,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b111001; i1 = 6'b010111; // Expected: {'sum': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b111001; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 3101,
                 
                 sum
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b011111; i1 = 6'b011011; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b011111; i1 = 6'b011011; | Outputs: sum=%b | Expected: sum=%d",
                 3102,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b110101; i1 = 6'b110101; // Expected: {'sum': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b110101; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 3103,
                 
                 sum
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b110101; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b110101; | Outputs: sum=%b | Expected: sum=%d",
                 3104,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b100011; i1 = 6'b101010; // Expected: {'sum': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b100011; i1 = 6'b101010; | Outputs: sum=%b | Expected: sum=%d",
                 3105,
                 
                 sum
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100100; i1 = 6'b001001; // Expected: {'sum': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100100; i1 = 6'b001001; | Outputs: sum=%b | Expected: sum=%d",
                 3106,
                 
                 sum
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b101101; // Expected: {'sum': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 3107,
                 
                 sum
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010101; i1 = 6'b100101; // Expected: {'sum': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010101; i1 = 6'b100101; | Outputs: sum=%b | Expected: sum=%d",
                 3108,
                 
                 sum
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b001110; i1 = 6'b110100; // Expected: {'sum': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b001110; i1 = 6'b110100; | Outputs: sum=%b | Expected: sum=%d",
                 3109,
                 
                 sum
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001001; i1 = 6'b000101; // Expected: {'sum': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001001; i1 = 6'b000101; | Outputs: sum=%b | Expected: sum=%d",
                 3110,
                 
                 sum
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b110010; i1 = 6'b110110; // Expected: {'sum': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b110010; i1 = 6'b110110; | Outputs: sum=%b | Expected: sum=%d",
                 3111,
                 
                 sum
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b011110; i1 = 6'b000110; // Expected: {'sum': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b011110; i1 = 6'b000110; | Outputs: sum=%b | Expected: sum=%d",
                 3112,
                 
                 sum
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b101011; i1 = 6'b101101; // Expected: {'sum': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b101011; i1 = 6'b101101; | Outputs: sum=%b | Expected: sum=%d",
                 3113,
                 
                 sum
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100011; i1 = 6'b000111; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100011; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 3114,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010010; i1 = 6'b001100; // Expected: {'sum': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010010; i1 = 6'b001100; | Outputs: sum=%b | Expected: sum=%d",
                 3115,
                 
                 sum
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b010110; i1 = 6'b101001; // Expected: {'sum': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b010110; i1 = 6'b101001; | Outputs: sum=%b | Expected: sum=%d",
                 3116,
                 
                 sum
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b100011; i1 = 6'b010111; // Expected: {'sum': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b100011; i1 = 6'b010111; | Outputs: sum=%b | Expected: sum=%d",
                 3117,
                 
                 sum
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b101001; i1 = 6'b001101; // Expected: {'sum': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b101001; i1 = 6'b001101; | Outputs: sum=%b | Expected: sum=%d",
                 3118,
                 
                 sum
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010000; i1 = 6'b100011; // Expected: {'sum': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010000; i1 = 6'b100011; | Outputs: sum=%b | Expected: sum=%d",
                 3119,
                 
                 sum
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b1; i0 = 6'b001111; i1 = 6'b000111; // Expected: {'sum': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b1; i0 = 6'b001111; i1 = 6'b000111; | Outputs: sum=%b | Expected: sum=%d",
                 3120,
                 
                 sum
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 cin = 1'b0; i0 = 6'b010111; i1 = 6'b011111; // Expected: {'sum': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: cin = 1'b0; i0 = 6'b010111; i1 = 6'b011111; | Outputs: sum=%b | Expected: sum=%d",
                 3121,
                 
                 sum
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        $finish;
    end
  
endmodule