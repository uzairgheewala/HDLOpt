
`timescale 1ns / 1ps

module tb_N8_booth_multiplier;

    // Parameters
    
    parameter N = 8;
    
     
    // Inputs
    
    reg   clk;
    
    reg   rst;
    
    reg   start;
    
    reg signed [7:0] X;
    
    reg signed [7:0] Y;
    
    
    // Outputs
    
    wire signed [15:0] Z;
    
    wire   valid;
    
    
    // Instantiate the Unit Under Test (UUT)
    booth_multiplier  #( N ) uut (
        
        .clk(clk),
        
        .rst(rst),
        
        .start(start),
        
        .X(X),
        
        .Y(Y),
        
        
        .Z(Z),
        
        .valid(valid)
        
    );

    // Clock generation 
    
    
            always begin
                #5 clk = ~clk;
            end
            
    

    
    
            always begin
                #99 rst = 1'b1; 
            end
            
    
    
    initial begin
        // Initialize Inputs
        
        clk = 0;
        
        rst = 0;
        
        start = 0;
        
        X = 0;
        
        Y = 0;
        
    
        // Wait for global reset
        #100;
    
        // Stimuli
        
        #10 X = 8'b11011010; Y = 8'b01000000; // Expected: {'Z': -2432}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011010; Y = 8'b01000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 0,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001110; Y = 8'b01001000; // Expected: {'Z': -3600}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001110; Y = 8'b01001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011001; Y = 8'b11010110; // Expected: {'Z': 4326}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011001; Y = 8'b11010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4326
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001100; Y = 8'b11100010; // Expected: {'Z': 3480}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001100; Y = 8'b11100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000100; Y = 8'b10010011; // Expected: {'Z': -436}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000100; Y = 8'b10010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 4,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -436
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b10101010; // Expected: {'Z': -1118}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b10101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 5,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110000; Y = 8'b00011101; // Expected: {'Z': -464}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110000; Y = 8'b00011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 6,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111011; Y = 8'b10100110; // Expected: {'Z': -5310}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111011; Y = 8'b10100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 7,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5310
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001111; Y = 8'b00010010; // Expected: {'Z': -2034}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001111; Y = 8'b00010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 8,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2034
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b10101100; // Expected: {'Z': -3276}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b10101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 9,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3276
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110011; Y = 8'b11000110; // Expected: {'Z': -6670}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110011; Y = 8'b11000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 10,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6670
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b11011100; // Expected: {'Z': -1944}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b11011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 11,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010000; Y = 8'b10110001; // Expected: {'Z': 3792}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010000; Y = 8'b10110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 12,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001010; Y = 8'b01111100; // Expected: {'Z': -6696}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001010; Y = 8'b01111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 13,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6696
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110111; Y = 8'b01001100; // Expected: {'Z': -684}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110111; Y = 8'b01001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 14,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -684
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100011; Y = 8'b11101000; // Expected: {'Z': -2376}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100011; Y = 8'b11101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 15,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2376
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b10001000; // Expected: {'Z': -6480}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b10001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 16,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011110; Y = 8'b10101111; // Expected: {'Z': -2430}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011110; Y = 8'b10101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 17,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001100; Y = 8'b10100010; // Expected: {'Z': 10904}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001100; Y = 8'b10100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 18,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10904
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001011; Y = 8'b00001001; // Expected: {'Z': -1053}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001011; Y = 8'b00001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 19,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1053
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100101; Y = 8'b00110000; // Expected: {'Z': 1776}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100101; Y = 8'b00110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 20,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1776
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011111; Y = 8'b10011101; // Expected: {'Z': 9603}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011111; Y = 8'b10011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 21,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9603
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111011; Y = 8'b10000000; // Expected: {'Z': -7552}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111011; Y = 8'b10000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 22,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b10111001; // Expected: {'Z': -4828}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b10111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 23,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011011; Y = 8'b01011010; // Expected: {'Z': 8190}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011011; Y = 8'b01011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 24,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001001; Y = 8'b11011100; // Expected: {'Z': -2628}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001001; Y = 8'b11011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 25,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2628
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110101; Y = 8'b10100111; // Expected: {'Z': 979}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110101; Y = 8'b10100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 26,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 979
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111001; Y = 8'b00011010; // Expected: {'Z': -182}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111001; Y = 8'b00011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 27,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000000; Y = 8'b00101010; // Expected: {'Z': -5376}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000000; Y = 8'b00101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 28,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5376
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000111; Y = 8'b10100100; // Expected: {'Z': -644}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000111; Y = 8'b10100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 29,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -644
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111000; Y = 8'b10111001; // Expected: {'Z': -8520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111000; Y = 8'b10111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 30,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111110; Y = 8'b10110001; // Expected: {'Z': 5214}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111110; Y = 8'b10110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 31,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011001; Y = 8'b11110111; // Expected: {'Z': -225}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011001; Y = 8'b11110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 32,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001011; Y = 8'b01001110; // Expected: {'Z': -4134}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001011; Y = 8'b01001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 33,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b10101111; // Expected: {'Z': -7128}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b10101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 34,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b11010000; // Expected: {'Z': -912}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b11010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 35,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -912
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010101; Y = 8'b10101101; // Expected: {'Z': -7055}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010101; Y = 8'b10101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 36,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7055
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001101; Y = 8'b11010111; // Expected: {'Z': -3157}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001101; Y = 8'b11010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 37,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3157
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001111; Y = 8'b00011010; // Expected: {'Z': -1274}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001111; Y = 8'b00011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 38,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1274
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101000; Y = 8'b00001001; // Expected: {'Z': 360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101000; Y = 8'b00001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 39,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011011; Y = 8'b01011101; // Expected: {'Z': -9393}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011011; Y = 8'b01011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 40,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9393
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011101; Y = 8'b11110101; // Expected: {'Z': 385}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011101; Y = 8'b11110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 41,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 385
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000100; Y = 8'b10101011; // Expected: {'Z': 5100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000100; Y = 8'b10101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 42,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b11111101; // Expected: {'Z': -39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b11111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 43,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b01010110; // Expected: {'Z': -9546}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b01010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 44,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011110; Y = 8'b11101100; // Expected: {'Z': -1880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011110; Y = 8'b11101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 45,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100100; Y = 8'b01000111; // Expected: {'Z': 7100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100100; Y = 8'b01000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 46,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110110; Y = 8'b11100000; // Expected: {'Z': 2368}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110110; Y = 8'b11100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 47,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001101; Y = 8'b11010011; // Expected: {'Z': 5175}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001101; Y = 8'b11010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 48,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100101; Y = 8'b00011101; // Expected: {'Z': 2929}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100101; Y = 8'b00011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 49,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2929
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100101; Y = 8'b11111101; // Expected: {'Z': 273}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100101; Y = 8'b11111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 50,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 273
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110100; Y = 8'b00100101; // Expected: {'Z': 4292}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110100; Y = 8'b00100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 51,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4292
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100010; Y = 8'b10111101; // Expected: {'Z': -6566}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100010; Y = 8'b10111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 52,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6566
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011110; Y = 8'b00101011; // Expected: {'Z': -1462}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011110; Y = 8'b00101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 53,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110100; Y = 8'b01110010; // Expected: {'Z': -1368}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110100; Y = 8'b01110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 54,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b00000110; // Expected: {'Z': -354}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b00000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 55,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -354
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111111; Y = 8'b10101101; // Expected: {'Z': 83}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111111; Y = 8'b10101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 56,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011111; Y = 8'b11101000; // Expected: {'Z': -2280}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011111; Y = 8'b11101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 57,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011101; Y = 8'b11110000; // Expected: {'Z': 1584}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011101; Y = 8'b11110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 58,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1584
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011110; Y = 8'b11000011; // Expected: {'Z': 5978}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011110; Y = 8'b11000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 59,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5978
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010110; Y = 8'b10101010; // Expected: {'Z': -7396}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010110; Y = 8'b10101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 60,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7396
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011000; Y = 8'b11000011; // Expected: {'Z': 2440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011000; Y = 8'b11000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 61,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011100; Y = 8'b00101101; // Expected: {'Z': 1260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011100; Y = 8'b00101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 62,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010000; Y = 8'b00011011; // Expected: {'Z': -3024}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010000; Y = 8'b00011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 63,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010101; Y = 8'b00011010; // Expected: {'Z': 2210}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010101; Y = 8'b00011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 64,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100011; Y = 8'b11011110; // Expected: {'Z': -3366}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100011; Y = 8'b11011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 65,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3366
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001111; Y = 8'b01001011; // Expected: {'Z': -3675}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001111; Y = 8'b01001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 66,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3675
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100110; Y = 8'b11110100; // Expected: {'Z': 1080}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100110; Y = 8'b11110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 67,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b01111001; // Expected: {'Z': -10164}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b01111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 68,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101011; Y = 8'b00101010; // Expected: {'Z': -3570}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101011; Y = 8'b00101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 69,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3570
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101111; Y = 8'b01011110; // Expected: {'Z': 10434}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101111; Y = 8'b01011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 70,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10434
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100000; Y = 8'b00110011; // Expected: {'Z': -4896}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100000; Y = 8'b00110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 71,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b01110010; // Expected: {'Z': 10032}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b01110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 72,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10032
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011011; Y = 8'b11001110; // Expected: {'Z': -1350}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011011; Y = 8'b11001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 73,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110001; Y = 8'b00110110; // Expected: {'Z': 2646}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110001; Y = 8'b00110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 74,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2646
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001000; Y = 8'b00100010; // Expected: {'Z': 272}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001000; Y = 8'b00100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 75,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 272
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011000; Y = 8'b10111011; // Expected: {'Z': -1656}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011000; Y = 8'b10111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 76,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1656
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000011; Y = 8'b10101100; // Expected: {'Z': 10500}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000011; Y = 8'b10101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 77,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011010; Y = 8'b11110110; // Expected: {'Z': 1020}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011010; Y = 8'b11110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 78,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1020
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110111; Y = 8'b11011000; // Expected: {'Z': 2920}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110111; Y = 8'b11011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 79,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001110; Y = 8'b01000101; // Expected: {'Z': 966}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001110; Y = 8'b01000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 80,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 966
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000010; Y = 8'b00111010; // Expected: {'Z': -3596}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000010; Y = 8'b00111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 81,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3596
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110000; Y = 8'b00000010; // Expected: {'Z': -160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110000; Y = 8'b00000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 82,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010110; Y = 8'b10011101; // Expected: {'Z': 4158}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010110; Y = 8'b10011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 83,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4158
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100011; Y = 8'b11010111; // Expected: {'Z': 1189}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100011; Y = 8'b11010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 84,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001110; Y = 8'b11111100; // Expected: {'Z': -56}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001110; Y = 8'b11111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 85,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011100; Y = 8'b11110010; // Expected: {'Z': -1288}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011100; Y = 8'b11110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 86,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111100; Y = 8'b01101010; // Expected: {'Z': 13144}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111100; Y = 8'b01101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 87,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 13144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101110; Y = 8'b10010000; // Expected: {'Z': -5152}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101110; Y = 8'b10010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 88,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b00010110; // Expected: {'Z': -1232}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b00010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 89,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001100; Y = 8'b10011100; // Expected: {'Z': 5200}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001100; Y = 8'b10011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 90,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001010; Y = 8'b10011001; // Expected: {'Z': -1030}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001010; Y = 8'b10011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 91,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1030
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b01110110; // Expected: {'Z': 7198}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b01110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 92,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000010; Y = 8'b01111111; // Expected: {'Z': -16002}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000010; Y = 8'b01111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 93,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -16002
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b10000000; // Expected: {'Z': -2432}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b10000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 94,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011010; Y = 8'b10101111; // Expected: {'Z': 8262}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011010; Y = 8'b10101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 95,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8262
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b11011011; // Expected: {'Z': -2516}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b11011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 96,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2516
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011011; Y = 8'b10001100; // Expected: {'Z': -3132}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011011; Y = 8'b10001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 97,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001110; Y = 8'b11101101; // Expected: {'Z': -266}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001110; Y = 8'b11101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 98,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -266
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b01001010; // Expected: {'Z': -6068}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b01001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 99,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6068
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111100; Y = 8'b10001101; // Expected: {'Z': 460}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111100; Y = 8'b10001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 100,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 460
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b00100110; // Expected: {'Z': 4674}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b00100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 101,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4674
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101011; Y = 8'b01111101; // Expected: {'Z': 5375}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101011; Y = 8'b01111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 102,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5375
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110001; Y = 8'b00111001; // Expected: {'Z': -855}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110001; Y = 8'b00111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 103,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -855
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111110; Y = 8'b10010001; // Expected: {'Z': 222}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111110; Y = 8'b10010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 104,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b00010111; // Expected: {'Z': 2208}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b00010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 105,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110100; Y = 8'b11001100; // Expected: {'Z': 3952}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110100; Y = 8'b11001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 106,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3952
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001101; Y = 8'b10010010; // Expected: {'Z': -8470}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001101; Y = 8'b10010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 107,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8470
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100110; Y = 8'b10100000; // Expected: {'Z': 8640}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100110; Y = 8'b10100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 108,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100101; Y = 8'b00110000; // Expected: {'Z': -4368}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100101; Y = 8'b00110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 109,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110110; Y = 8'b10101100; // Expected: {'Z': 840}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110110; Y = 8'b10101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 110,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110000; Y = 8'b10011001; // Expected: {'Z': 8240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110000; Y = 8'b10011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 111,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b11000101; // Expected: {'Z': -3186}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b11000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 112,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111000; Y = 8'b00000010; // Expected: {'Z': 112}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111000; Y = 8'b00000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 113,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100101; Y = 8'b00011101; // Expected: {'Z': 1073}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100101; Y = 8'b00011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 114,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1073
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100010; Y = 8'b01100011; // Expected: {'Z': 3366}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100010; Y = 8'b01100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 115,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3366
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110011; Y = 8'b00011101; // Expected: {'Z': 3335}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110011; Y = 8'b00011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 116,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3335
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111010; Y = 8'b10101010; // Expected: {'Z': 516}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111010; Y = 8'b10101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 117,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 516
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000001; Y = 8'b01010010; // Expected: {'Z': -5166}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000001; Y = 8'b01010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 118,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100001; Y = 8'b01101001; // Expected: {'Z': 10185}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100001; Y = 8'b01101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 119,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111000; Y = 8'b00000110; // Expected: {'Z': -432}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111000; Y = 8'b00000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 120,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101010; Y = 8'b01100110; // Expected: {'Z': 4284}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101010; Y = 8'b01100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 121,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4284
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110111; Y = 8'b00010111; // Expected: {'Z': -1679}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110111; Y = 8'b00010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 122,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1679
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101110; Y = 8'b01110011; // Expected: {'Z': 5290}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101110; Y = 8'b01110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 123,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5290
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111010; Y = 8'b10010110; // Expected: {'Z': 7420}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111010; Y = 8'b10010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 124,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b10001011; // Expected: {'Z': 7956}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b10001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 125,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7956
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000010; Y = 8'b11011001; // Expected: {'Z': -2574}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000010; Y = 8'b11011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 126,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2574
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011001; Y = 8'b01100001; // Expected: {'Z': -9991}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011001; Y = 8'b01100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 127,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9991
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000100; Y = 8'b11001000; // Expected: {'Z': 6944}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000100; Y = 8'b11001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 128,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100110; Y = 8'b00001110; // Expected: {'Z': 1428}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100110; Y = 8'b00001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 129,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1428
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b00100100; // Expected: {'Z': 1692}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b00100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 130,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1692
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101011; Y = 8'b00100110; // Expected: {'Z': 4066}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101011; Y = 8'b00100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 131,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4066
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100010; Y = 8'b10000010; // Expected: {'Z': -12348}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100010; Y = 8'b10000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 132,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12348
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000010; Y = 8'b11110110; // Expected: {'Z': 620}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000010; Y = 8'b11110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 133,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110100; Y = 8'b10001010; // Expected: {'Z': -6136}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110100; Y = 8'b10001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 134,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111011; Y = 8'b00011110; // Expected: {'Z': -2070}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111011; Y = 8'b00011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 135,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2070
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100011; Y = 8'b01000000; // Expected: {'Z': 6336}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100011; Y = 8'b01000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 136,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6336
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100010; Y = 8'b10100100; // Expected: {'Z': -9016}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100010; Y = 8'b10100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 137,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b11010101; // Expected: {'Z': -2623}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b11010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 138,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2623
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000000; Y = 8'b10000101; // Expected: {'Z': 7872}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000000; Y = 8'b10000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 139,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7872
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100110; Y = 8'b00000001; // Expected: {'Z': -26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100110; Y = 8'b00000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 140,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100001; Y = 8'b00011011; // Expected: {'Z': 891}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100001; Y = 8'b00011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 141,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 891
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111111; Y = 8'b01011011; // Expected: {'Z': 11557}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111111; Y = 8'b01011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 142,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11557
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b10001001; // Expected: {'Z': -8092}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b10001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 143,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8092
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111100; Y = 8'b00101100; // Expected: {'Z': -176}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111100; Y = 8'b00101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 144,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111000; Y = 8'b01000110; // Expected: {'Z': 3920}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111000; Y = 8'b01000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 145,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001110; Y = 8'b10110010; // Expected: {'Z': 3900}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001110; Y = 8'b10110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 146,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100101; Y = 8'b01000111; // Expected: {'Z': 2627}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100101; Y = 8'b01000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 147,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2627
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011110; Y = 8'b10110010; // Expected: {'Z': -7332}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011110; Y = 8'b10110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 148,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7332
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011101; Y = 8'b11110000; // Expected: {'Z': 1584}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011101; Y = 8'b11110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 149,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1584
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101111; Y = 8'b00011011; // Expected: {'Z': 2997}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101111; Y = 8'b00011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 150,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2997
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101000; Y = 8'b11011110; // Expected: {'Z': -1360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101000; Y = 8'b11011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 151,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000011; Y = 8'b11111000; // Expected: {'Z': 488}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000011; Y = 8'b11111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 152,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110101; Y = 8'b01000000; // Expected: {'Z': 7488}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110101; Y = 8'b01000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 153,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111101; Y = 8'b01100001; // Expected: {'Z': -6499}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111101; Y = 8'b01100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 154,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6499
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101010; Y = 8'b01011100; // Expected: {'Z': -7912}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101010; Y = 8'b01011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 155,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7912
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110110; Y = 8'b00111100; // Expected: {'Z': -4440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110110; Y = 8'b00111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 156,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100101; Y = 8'b00101010; // Expected: {'Z': 1554}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100101; Y = 8'b00101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 157,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1554
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110100; Y = 8'b10111101; // Expected: {'Z': -7772}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110100; Y = 8'b10111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 158,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7772
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b00010110; // Expected: {'Z': 792}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b00010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 159,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110001; Y = 8'b10000101; // Expected: {'Z': 1845}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110001; Y = 8'b10000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 160,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1845
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101011; Y = 8'b10110011; // Expected: {'Z': 1617}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101011; Y = 8'b10110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 161,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1617
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100011; Y = 8'b11000011; // Expected: {'Z': 5673}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100011; Y = 8'b11000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 162,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5673
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011101; Y = 8'b11000110; // Expected: {'Z': 2030}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011101; Y = 8'b11000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 163,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2030
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001101; Y = 8'b11101101; // Expected: {'Z': -1463}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001101; Y = 8'b11101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 164,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1463
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111000; Y = 8'b10011010; // Expected: {'Z': -12240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111000; Y = 8'b10011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 165,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100001; Y = 8'b00111010; // Expected: {'Z': 5626}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100001; Y = 8'b00111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 166,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5626
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011100; Y = 8'b10100101; // Expected: {'Z': -8372}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011100; Y = 8'b10100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 167,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8372
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101110; Y = 8'b01100011; // Expected: {'Z': -1782}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101110; Y = 8'b01100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 168,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1782
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111001; Y = 8'b00101111; // Expected: {'Z': 5687}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111001; Y = 8'b00101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 169,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5687
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001111; Y = 8'b00011011; // Expected: {'Z': -1323}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001111; Y = 8'b00011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 170,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1323
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000101; Y = 8'b11010010; // Expected: {'Z': -230}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000101; Y = 8'b11010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 171,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000110; Y = 8'b01010100; // Expected: {'Z': -4872}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000110; Y = 8'b01010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 172,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4872
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b00100111; // Expected: {'Z': -3276}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b00100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 173,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3276
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000100; Y = 8'b01001100; // Expected: {'Z': -4560}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000100; Y = 8'b01001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 174,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110101; Y = 8'b11001011; // Expected: {'Z': -2809}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110101; Y = 8'b11001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 175,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2809
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011100; Y = 8'b10011001; // Expected: {'Z': -2884}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011100; Y = 8'b10011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 176,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2884
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001010; Y = 8'b01110111; // Expected: {'Z': -6426}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001010; Y = 8'b01110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 177,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6426
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001011; Y = 8'b00110101; // Expected: {'Z': -2809}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001011; Y = 8'b00110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 178,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2809
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001010; Y = 8'b10001100; // Expected: {'Z': 13688}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001010; Y = 8'b10001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 179,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 13688
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111000; Y = 8'b10001010; // Expected: {'Z': 944}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111000; Y = 8'b10001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 180,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b11000000; // Expected: {'Z': 3584}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b11000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 181,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3584
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011111; Y = 8'b11011111; // Expected: {'Z': -3135}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011111; Y = 8'b11011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 182,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000010; Y = 8'b10000100; // Expected: {'Z': -8184}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000010; Y = 8'b10000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 183,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110100; Y = 8'b00000111; // Expected: {'Z': -532}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110100; Y = 8'b00000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 184,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -532
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001100; Y = 8'b10001000; // Expected: {'Z': -1440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001100; Y = 8'b10001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 185,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000001; Y = 8'b11101000; // Expected: {'Z': 3048}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000001; Y = 8'b11101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 186,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3048
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011000; Y = 8'b00010001; // Expected: {'Z': 408}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011000; Y = 8'b00010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 187,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110001; Y = 8'b11100010; // Expected: {'Z': 2370}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110001; Y = 8'b11100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 188,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2370
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100101; Y = 8'b11101100; // Expected: {'Z': -2020}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100101; Y = 8'b11101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 189,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2020
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111000; Y = 8'b10011000; // Expected: {'Z': 7488}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111000; Y = 8'b10011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 190,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011110; Y = 8'b10101100; // Expected: {'Z': 2856}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011110; Y = 8'b10101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 191,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110010; Y = 8'b00011111; // Expected: {'Z': 3534}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110010; Y = 8'b00011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 192,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3534
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b10100110; // Expected: {'Z': -11070}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b10100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 193,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11070
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010010; Y = 8'b01001100; // Expected: {'Z': 1368}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010010; Y = 8'b01001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 194,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110111; Y = 8'b11100010; // Expected: {'Z': -1650}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110111; Y = 8'b11100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 195,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100101; Y = 8'b01101100; // Expected: {'Z': -9828}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100101; Y = 8'b01101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 196,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b10100001; // Expected: {'Z': -2755}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b10100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 197,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2755
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100001; Y = 8'b01010110; // Expected: {'Z': -8170}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100001; Y = 8'b01010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 198,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100111; Y = 8'b01101010; // Expected: {'Z': -9434}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100111; Y = 8'b01101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 199,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9434
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000000; Y = 8'b00010011; // Expected: {'Z': -2432}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000000; Y = 8'b00010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 200,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001001; Y = 8'b10111011; // Expected: {'Z': -5037}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001001; Y = 8'b10111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 201,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5037
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111100; Y = 8'b10101000; // Expected: {'Z': -5280}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111100; Y = 8'b10101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 202,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011011; Y = 8'b01011001; // Expected: {'Z': 8099}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011011; Y = 8'b01011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 203,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8099
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001111; Y = 8'b10000000; // Expected: {'Z': 6272}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001111; Y = 8'b10000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 204,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6272
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000110; Y = 8'b10111000; // Expected: {'Z': -5040}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000110; Y = 8'b10111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 205,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111111; Y = 8'b10010101; // Expected: {'Z': 107}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111111; Y = 8'b10010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 206,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110110; Y = 8'b00111011; // Expected: {'Z': -590}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110110; Y = 8'b00111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 207,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -590
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111001; Y = 8'b10111110; // Expected: {'Z': -7986}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111001; Y = 8'b10111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 208,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7986
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001110; Y = 8'b01101110; // Expected: {'Z': -12540}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001110; Y = 8'b01101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 209,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b00101110; // Expected: {'Z': 3128}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b00101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 210,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101010; Y = 8'b00010111; // Expected: {'Z': 2438}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101010; Y = 8'b00010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 211,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2438
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111101; Y = 8'b00110001; // Expected: {'Z': -147}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111101; Y = 8'b00110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 212,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010101; Y = 8'b01011000; // Expected: {'Z': -9416}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010101; Y = 8'b01011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 213,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101011; Y = 8'b00011010; // Expected: {'Z': -546}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101011; Y = 8'b00011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 214,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100110; Y = 8'b10001011; // Expected: {'Z': -11934}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100110; Y = 8'b10001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 215,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11934
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011111; Y = 8'b00000011; // Expected: {'Z': 93}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011111; Y = 8'b00000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 216,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001111; Y = 8'b10000101; // Expected: {'Z': 13899}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001111; Y = 8'b10000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 217,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 13899
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001101; Y = 8'b11000111; // Expected: {'Z': -4389}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001101; Y = 8'b11000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 218,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4389
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000100; Y = 8'b11111101; // Expected: {'Z': 372}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000100; Y = 8'b11111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 219,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 372
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001111; Y = 8'b01000100; // Expected: {'Z': -7684}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001111; Y = 8'b01000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 220,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7684
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010111; Y = 8'b11111000; // Expected: {'Z': -696}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010111; Y = 8'b11111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 221,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -696
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010111; Y = 8'b10110000; // Expected: {'Z': -1840}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010111; Y = 8'b10110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 222,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110111; Y = 8'b10100100; // Expected: {'Z': -5060}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110111; Y = 8'b10100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 223,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000110; Y = 8'b01110011; // Expected: {'Z': 8050}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000110; Y = 8'b01110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 224,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000100; Y = 8'b01111111; // Expected: {'Z': -7620}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000100; Y = 8'b01111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 225,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100001; Y = 8'b00101110; // Expected: {'Z': -4370}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100001; Y = 8'b00101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 226,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4370
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110111; Y = 8'b00000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110111; Y = 8'b00000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 227,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100011; Y = 8'b00101000; // Expected: {'Z': -1160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100011; Y = 8'b00101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 228,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b10101101; // Expected: {'Z': -8549}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b10101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 229,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8549
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100111; Y = 8'b11110011; // Expected: {'Z': 325}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100111; Y = 8'b11110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 230,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 325
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111111; Y = 8'b10011100; // Expected: {'Z': -6300}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111111; Y = 8'b10011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 231,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010100; Y = 8'b00000011; // Expected: {'Z': -324}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010100; Y = 8'b00000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 232,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -324
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110011; Y = 8'b01111000; // Expected: {'Z': 6120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110011; Y = 8'b01111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 233,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110111; Y = 8'b01110100; // Expected: {'Z': -8468}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110111; Y = 8'b01110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 234,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8468
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110011; Y = 8'b10111111; // Expected: {'Z': 5005}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110011; Y = 8'b10111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 235,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5005
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100001; Y = 8'b11011011; // Expected: {'Z': -1221}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100001; Y = 8'b11011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 236,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001011; Y = 8'b10110011; // Expected: {'Z': -5775}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001011; Y = 8'b10110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 237,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5775
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010101; Y = 8'b00011011; // Expected: {'Z': -2889}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010101; Y = 8'b00011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 238,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2889
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b00100100; // Expected: {'Z': -2952}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b00100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 239,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2952
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011010; Y = 8'b11011011; // Expected: {'Z': 3774}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011010; Y = 8'b11011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 240,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3774
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110101; Y = 8'b11100110; // Expected: {'Z': -1378}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110101; Y = 8'b11100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 241,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1378
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b00111100; // Expected: {'Z': 1140}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b00111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 242,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110101; Y = 8'b00011110; // Expected: {'Z': -330}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110101; Y = 8'b00011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 243,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -330
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000101; Y = 8'b00100001; // Expected: {'Z': 165}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000101; Y = 8'b00100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 244,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111110; Y = 8'b00011010; // Expected: {'Z': 3276}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111110; Y = 8'b00011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 245,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3276
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101000; Y = 8'b11001011; // Expected: {'Z': -2120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101000; Y = 8'b11001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 246,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110001; Y = 8'b00110101; // Expected: {'Z': -795}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110001; Y = 8'b00110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 247,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -795
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100010; Y = 8'b00011010; // Expected: {'Z': 884}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100010; Y = 8'b00011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 248,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 884
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000000; Y = 8'b10010000; // Expected: {'Z': 7168}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000000; Y = 8'b10010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 249,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110111; Y = 8'b01001010; // Expected: {'Z': 8806}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110111; Y = 8'b01001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 250,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8806
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001100; Y = 8'b10001101; // Expected: {'Z': -1380}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001100; Y = 8'b10001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 251,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1380
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010010; Y = 8'b10000001; // Expected: {'Z': 13970}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010010; Y = 8'b10000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 252,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 13970
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100001; Y = 8'b10001010; // Expected: {'Z': 3658}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100001; Y = 8'b10001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 253,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3658
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111111; Y = 8'b10110001; // Expected: {'Z': 79}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111111; Y = 8'b10110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 254,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101101; Y = 8'b00111110; // Expected: {'Z': 2790}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101101; Y = 8'b00111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 255,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2790
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011011; Y = 8'b00101111; // Expected: {'Z': 4277}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011011; Y = 8'b00101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 256,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4277
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000111; Y = 8'b00100110; // Expected: {'Z': 266}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000111; Y = 8'b00100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 257,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 266
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011110; Y = 8'b01101110; // Expected: {'Z': -10780}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011110; Y = 8'b01101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 258,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101011; Y = 8'b00101000; // Expected: {'Z': 1720}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101011; Y = 8'b00101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 259,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010011; Y = 8'b01110110; // Expected: {'Z': -5310}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010011; Y = 8'b01110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 260,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5310
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000100; Y = 8'b00010101; // Expected: {'Z': -2604}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000100; Y = 8'b00010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 261,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2604
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111001; Y = 8'b00100101; // Expected: {'Z': -2627}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111001; Y = 8'b00100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 262,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2627
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010100; Y = 8'b01100100; // Expected: {'Z': 2000}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010100; Y = 8'b01100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 263,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100110; Y = 8'b00010111; // Expected: {'Z': -2070}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100110; Y = 8'b00010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 264,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2070
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100101; Y = 8'b11110001; // Expected: {'Z': -555}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100101; Y = 8'b11110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 265,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -555
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110101; Y = 8'b00011011; // Expected: {'Z': -297}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110101; Y = 8'b00011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 266,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -297
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111001; Y = 8'b01011110; // Expected: {'Z': -658}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111001; Y = 8'b01011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 267,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -658
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b10011101; // Expected: {'Z': 10989}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b10011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 268,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10989
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101001; Y = 8'b01000011; // Expected: {'Z': 2747}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101001; Y = 8'b01000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 269,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2747
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000010; Y = 8'b10010110; // Expected: {'Z': 6572}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000010; Y = 8'b10010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 270,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6572
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010110; Y = 8'b00110011; // Expected: {'Z': 4386}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010110; Y = 8'b00110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 271,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4386
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111010; Y = 8'b10111101; // Expected: {'Z': -8174}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111010; Y = 8'b10111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 272,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010000; Y = 8'b11101101; // Expected: {'Z': -304}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010000; Y = 8'b11101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 273,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -304
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101001; Y = 8'b10011001; // Expected: {'Z': 2369}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101001; Y = 8'b10011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 274,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2369
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b01101101; // Expected: {'Z': 5123}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b01101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 275,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5123
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110001; Y = 8'b01100100; // Expected: {'Z': -7900}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110001; Y = 8'b01100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 276,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111010; Y = 8'b10010010; // Expected: {'Z': 660}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111010; Y = 8'b10010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 277,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110100; Y = 8'b00110101; // Expected: {'Z': 2756}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110100; Y = 8'b00110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 278,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001011; Y = 8'b00110100; // Expected: {'Z': 3900}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001011; Y = 8'b00110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 279,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110011; Y = 8'b01101000; // Expected: {'Z': -1352}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110011; Y = 8'b01101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 280,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001010; Y = 8'b00111101; // Expected: {'Z': 610}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001010; Y = 8'b00111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 281,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 610
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011010; Y = 8'b10001101; // Expected: {'Z': -2990}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011010; Y = 8'b10001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 282,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2990
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b01011011; // Expected: {'Z': 6188}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b01011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 283,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111001; Y = 8'b01111101; // Expected: {'Z': -8875}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111001; Y = 8'b01111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 284,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8875
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100001; Y = 8'b01100011; // Expected: {'Z': 9603}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100001; Y = 8'b01100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 285,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9603
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000010; Y = 8'b10000110; // Expected: {'Z': 7564}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000010; Y = 8'b10000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 286,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7564
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b00011111; // Expected: {'Z': -3441}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b00011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 287,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3441
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001101; Y = 8'b10010100; // Expected: {'Z': -8316}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001101; Y = 8'b10010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 288,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8316
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111101; Y = 8'b00101011; // Expected: {'Z': -2881}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111101; Y = 8'b00101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 289,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2881
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111010; Y = 8'b10011011; // Expected: {'Z': 7070}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111010; Y = 8'b10011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 290,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7070
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111001; Y = 8'b00101001; // Expected: {'Z': -287}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111001; Y = 8'b00101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 291,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -287
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000010; Y = 8'b11010110; // Expected: {'Z': 5292}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000010; Y = 8'b11010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 292,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5292
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010101; Y = 8'b00101010; // Expected: {'Z': -1806}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010101; Y = 8'b00101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 293,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1806
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011011; Y = 8'b11101111; // Expected: {'Z': -1547}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011011; Y = 8'b11101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 294,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1547
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000111; Y = 8'b01111111; // Expected: {'Z': -15367}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000111; Y = 8'b01111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 295,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -15367
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000110; Y = 8'b00010101; // Expected: {'Z': -1218}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000110; Y = 8'b00010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 296,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010101; Y = 8'b10111000; // Expected: {'Z': 7704}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010101; Y = 8'b10111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 297,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7704
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100101; Y = 8'b10001100; // Expected: {'Z': 3132}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100101; Y = 8'b10001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 298,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111111; Y = 8'b10101000; // Expected: {'Z': 88}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111111; Y = 8'b10101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 299,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b01010011; // Expected: {'Z': 3237}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b01010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 300,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3237
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100011; Y = 8'b01010111; // Expected: {'Z': 3045}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100011; Y = 8'b01010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 301,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3045
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110011; Y = 8'b11010010; // Expected: {'Z': 3542}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110011; Y = 8'b11010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 302,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3542
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010110; Y = 8'b01101011; // Expected: {'Z': -4494}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010110; Y = 8'b01101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 303,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4494
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011000; Y = 8'b11011001; // Expected: {'Z': 4056}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011000; Y = 8'b11011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 304,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4056
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001110; Y = 8'b11011010; // Expected: {'Z': -532}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001110; Y = 8'b11011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 305,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -532
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b11011111; // Expected: {'Z': -297}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b11011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 306,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -297
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111100; Y = 8'b00000011; // Expected: {'Z': 180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111100; Y = 8'b00000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 307,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000101; Y = 8'b01101001; // Expected: {'Z': 7245}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000101; Y = 8'b01101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 308,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011001; Y = 8'b11011000; // Expected: {'Z': 1560}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011001; Y = 8'b11011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 309,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110011; Y = 8'b01010011; // Expected: {'Z': -6391}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110011; Y = 8'b01010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 310,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6391
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011100; Y = 8'b00000010; // Expected: {'Z': 184}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011100; Y = 8'b00000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 311,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101000; Y = 8'b10100101; // Expected: {'Z': 8008}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101000; Y = 8'b10100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 312,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010101; Y = 8'b10010101; // Expected: {'Z': 4601}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010101; Y = 8'b10010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 313,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4601
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000001; Y = 8'b10001010; // Expected: {'Z': 7434}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000001; Y = 8'b10001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 314,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7434
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011110; Y = 8'b11011111; // Expected: {'Z': 3234}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011110; Y = 8'b11011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 315,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b10010111; // Expected: {'Z': -3780}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b10010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 316,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100101; Y = 8'b01010110; // Expected: {'Z': 8686}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100101; Y = 8'b01010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 317,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8686
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001110; Y = 8'b01101000; // Expected: {'Z': -11856}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001110; Y = 8'b01101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 318,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b11110111; // Expected: {'Z': -81}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b11110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 319,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000110; Y = 8'b11010011; // Expected: {'Z': 5490}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000110; Y = 8'b11010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 320,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5490
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111101; Y = 8'b00011000; // Expected: {'Z': -1608}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111101; Y = 8'b00011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 321,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1608
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001010; Y = 8'b01110110; // Expected: {'Z': -13924}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001010; Y = 8'b01110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 322,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -13924
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100101; Y = 8'b01010101; // Expected: {'Z': -2295}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100101; Y = 8'b01010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 323,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2295
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000111; Y = 8'b00001001; // Expected: {'Z': -1089}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000111; Y = 8'b00001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 324,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1089
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101110; Y = 8'b11011100; // Expected: {'Z': -1656}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101110; Y = 8'b11011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 325,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1656
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b01111001; // Expected: {'Z': 12463}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b01111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 326,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 12463
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b01101101; // Expected: {'Z': 218}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b01101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 327,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110100; Y = 8'b11011010; // Expected: {'Z': -4408}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110100; Y = 8'b11011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 328,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b00100101; // Expected: {'Z': -4107}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b00100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 329,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011101; Y = 8'b01110000; // Expected: {'Z': -11088}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011101; Y = 8'b01110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 330,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11088
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000010; Y = 8'b00010001; // Expected: {'Z': -1054}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000010; Y = 8'b00010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 331,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1054
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101001; Y = 8'b11001001; // Expected: {'Z': -2255}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101001; Y = 8'b11001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 332,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001100; Y = 8'b10011011; // Expected: {'Z': -1212}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001100; Y = 8'b10011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 333,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101011; Y = 8'b00111100; // Expected: {'Z': 6420}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101011; Y = 8'b00111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 334,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000111; Y = 8'b10011101; // Expected: {'Z': 11979}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000111; Y = 8'b10011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 335,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11979
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010011; Y = 8'b11110011; // Expected: {'Z': 1417}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010011; Y = 8'b11110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 336,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1417
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101011; Y = 8'b01001000; // Expected: {'Z': -1512}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101011; Y = 8'b01001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 337,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1512
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000111; Y = 8'b10001101; // Expected: {'Z': 13915}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000111; Y = 8'b10001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 338,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 13915
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000101; Y = 8'b11111010; // Expected: {'Z': -30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000101; Y = 8'b11111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 339,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b10100110; // Expected: {'Z': -180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b10100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 340,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001001; Y = 8'b10010010; // Expected: {'Z': 6050}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001001; Y = 8'b10010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 341,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b00111111; // Expected: {'Z': -5166}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b00111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 342,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000010; Y = 8'b10100101; // Expected: {'Z': 11466}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000010; Y = 8'b10100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 343,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11466
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010011; Y = 8'b00000111; // Expected: {'Z': -315}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010011; Y = 8'b00000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 344,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -315
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110011; Y = 8'b00111111; // Expected: {'Z': 3213}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110011; Y = 8'b00111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 345,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b11000111; // Expected: {'Z': 4674}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b11000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 346,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4674
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110001; Y = 8'b01011000; // Expected: {'Z': 4312}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110001; Y = 8'b01011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 347,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4312
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111001; Y = 8'b11000101; // Expected: {'Z': -3363}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111001; Y = 8'b11000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 348,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3363
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110010; Y = 8'b11110110; // Expected: {'Z': 780}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110010; Y = 8'b11110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 349,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010011; Y = 8'b01010011; // Expected: {'Z': 6889}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010011; Y = 8'b01010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 350,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6889
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111010; Y = 8'b10001101; // Expected: {'Z': 8050}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111010; Y = 8'b10001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 351,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110100; Y = 8'b00011011; // Expected: {'Z': 3132}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110100; Y = 8'b00011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 352,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000110; Y = 8'b10101100; // Expected: {'Z': -5880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000110; Y = 8'b10101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 353,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000101; Y = 8'b11011011; // Expected: {'Z': 4551}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000101; Y = 8'b11011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 354,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4551
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001111; Y = 8'b01110000; // Expected: {'Z': 8848}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001111; Y = 8'b01110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 355,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101010; Y = 8'b01101110; // Expected: {'Z': -9460}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101010; Y = 8'b01101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 356,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9460
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100001; Y = 8'b11111011; // Expected: {'Z': 475}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100001; Y = 8'b11111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 357,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 475
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001100; Y = 8'b01000011; // Expected: {'Z': -3484}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001100; Y = 8'b01000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 358,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3484
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b10000110; // Expected: {'Z': 6832}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b10000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 359,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6832
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001111; Y = 8'b10111101; // Expected: {'Z': 3283}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001111; Y = 8'b10111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 360,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3283
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b10101011; // Expected: {'Z': -6120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b10101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 361,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b01000000; // Expected: {'Z': 3456}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b01000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 362,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010011; Y = 8'b11000101; // Expected: {'Z': -4897}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010011; Y = 8'b11000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 363,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4897
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101101; Y = 8'b00011001; // Expected: {'Z': 1125}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101101; Y = 8'b00011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 364,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010010; Y = 8'b10001001; // Expected: {'Z': 5474}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010010; Y = 8'b10001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 365,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5474
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110110; Y = 8'b01111101; // Expected: {'Z': -1250}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110110; Y = 8'b01111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 366,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b11010100; // Expected: {'Z': -3872}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b11010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 367,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3872
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b01100110; // Expected: {'Z': -8568}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b01100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 368,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8568
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111001; Y = 8'b10110110; // Expected: {'Z': -4218}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111001; Y = 8'b10110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 369,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111111; Y = 8'b11101111; // Expected: {'Z': -2159}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111111; Y = 8'b11101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 370,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b10110000; // Expected: {'Z': -3120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b10110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 371,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111010; Y = 8'b10101001; // Expected: {'Z': 6090}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111010; Y = 8'b10101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 372,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6090
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111110; Y = 8'b11111101; // Expected: {'Z': 198}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111110; Y = 8'b11111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 373,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101010; Y = 8'b11000100; // Expected: {'Z': -2520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101010; Y = 8'b11000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 374,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000110; Y = 8'b01100101; // Expected: {'Z': 7070}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000110; Y = 8'b01100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 375,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7070
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011000; Y = 8'b01011000; // Expected: {'Z': -3520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011000; Y = 8'b01011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 376,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110111; Y = 8'b10000100; // Expected: {'Z': 9052}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110111; Y = 8'b10000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 377,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9052
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b00111111; // Expected: {'Z': 4662}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b00111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 378,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4662
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010101; Y = 8'b00011101; // Expected: {'Z': -3103}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010101; Y = 8'b00011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 379,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011100; Y = 8'b11101000; // Expected: {'Z': 2400}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011100; Y = 8'b11101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 380,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101111; Y = 8'b10011101; // Expected: {'Z': 1683}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101111; Y = 8'b10011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 381,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1683
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011010; Y = 8'b11110000; // Expected: {'Z': -1440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011010; Y = 8'b11110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 382,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110010; Y = 8'b00100010; // Expected: {'Z': 3876}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110010; Y = 8'b00100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 383,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3876
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111110; Y = 8'b01000101; // Expected: {'Z': -138}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111110; Y = 8'b01000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 384,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100010; Y = 8'b01010100; // Expected: {'Z': -7896}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100010; Y = 8'b01010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 385,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110001; Y = 8'b11101100; // Expected: {'Z': 300}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110001; Y = 8'b11101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 386,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111111; Y = 8'b00001000; // Expected: {'Z': 1016}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111111; Y = 8'b00001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 387,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b01010000; // Expected: {'Z': 160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b01010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 388,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000101; Y = 8'b01001011; // Expected: {'Z': -9225}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000101; Y = 8'b01001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 389,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b10001001; // Expected: {'Z': -238}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b10001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 390,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111010; Y = 8'b11000110; // Expected: {'Z': -7076}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111010; Y = 8'b11000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 391,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7076
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b11010110; // Expected: {'Z': -1848}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b11010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 392,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001100; Y = 8'b00000001; // Expected: {'Z': 76}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001100; Y = 8'b00000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 393,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111110; Y = 8'b01000110; // Expected: {'Z': 4340}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111110; Y = 8'b01000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 394,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010001; Y = 8'b01100101; // Expected: {'Z': -4747}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010001; Y = 8'b01100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 395,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4747
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100110; Y = 8'b11010001; // Expected: {'Z': 1222}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100110; Y = 8'b11010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 396,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110110; Y = 8'b11010000; // Expected: {'Z': -5664}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110110; Y = 8'b11010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 397,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5664
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010000; Y = 8'b00001110; // Expected: {'Z': 224}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010000; Y = 8'b00001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 398,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011101; Y = 8'b01110000; // Expected: {'Z': -11088}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011101; Y = 8'b01110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 399,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11088
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100111; Y = 8'b10000100; // Expected: {'Z': 11036}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100111; Y = 8'b10000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 400,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11036
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100000; Y = 8'b10011010; // Expected: {'Z': 9792}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100000; Y = 8'b10011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 401,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011111; Y = 8'b11111110; // Expected: {'Z': 194}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011111; Y = 8'b11111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 402,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 194
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010010; Y = 8'b00111011; // Expected: {'Z': -6490}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010010; Y = 8'b00111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 403,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6490
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100111; Y = 8'b11111111; // Expected: {'Z': 89}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100111; Y = 8'b11111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 404,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 89
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100010; Y = 8'b11010110; // Expected: {'Z': -4116}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100010; Y = 8'b11010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 405,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111000; Y = 8'b01111110; // Expected: {'Z': -9072}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111000; Y = 8'b01111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 406,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9072
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b10001100; // Expected: {'Z': -10208}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b10001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 407,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101001; Y = 8'b00100000; // Expected: {'Z': 3360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101001; Y = 8'b00100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 408,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110011; Y = 8'b01110110; // Expected: {'Z': -1534}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110011; Y = 8'b01110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 409,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1534
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100111; Y = 8'b10101000; // Expected: {'Z': 2200}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100111; Y = 8'b10101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 410,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100101; Y = 8'b10010000; // Expected: {'Z': -4144}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100101; Y = 8'b10010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 411,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110101; Y = 8'b11001011; // Expected: {'Z': 583}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110101; Y = 8'b11001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 412,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 583
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001001; Y = 8'b10100111; // Expected: {'Z': 10591}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001001; Y = 8'b10100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 413,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10591
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111111; Y = 8'b00111101; // Expected: {'Z': 7747}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111111; Y = 8'b00111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 414,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7747
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000011; Y = 8'b11000110; // Expected: {'Z': 3538}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000011; Y = 8'b11000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 415,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3538
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110100; Y = 8'b10111011; // Expected: {'Z': -8004}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110100; Y = 8'b10111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 416,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8004
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b00111110; // Expected: {'Z': -5394}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b00111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 417,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5394
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001010; Y = 8'b11111000; // Expected: {'Z': -80}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001010; Y = 8'b11111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 418,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100011; Y = 8'b11111001; // Expected: {'Z': 651}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100011; Y = 8'b11111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 419,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 651
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011000; Y = 8'b10010100; // Expected: {'Z': -2592}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011000; Y = 8'b10010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 420,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2592
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b01111101; // Expected: {'Z': 8500}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b01111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 421,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010010; Y = 8'b00110110; // Expected: {'Z': -2484}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010010; Y = 8'b00110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 422,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2484
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111101; Y = 8'b10101000; // Expected: {'Z': 264}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111101; Y = 8'b10101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 423,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100101; Y = 8'b10010000; // Expected: {'Z': 3024}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100101; Y = 8'b10010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 424,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000111; Y = 8'b00100111; // Expected: {'Z': 2769}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000111; Y = 8'b00100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 425,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2769
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b11010010; // Expected: {'Z': -4416}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b11010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 426,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100011; Y = 8'b00000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100011; Y = 8'b00000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 427,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110001; Y = 8'b10001010; // Expected: {'Z': -13334}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110001; Y = 8'b10001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 428,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -13334
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110110; Y = 8'b10011001; // Expected: {'Z': 1030}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110110; Y = 8'b10011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 429,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1030
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001110; Y = 8'b00100000; // Expected: {'Z': -1600}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001110; Y = 8'b00100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 430,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011100; Y = 8'b10000101; // Expected: {'Z': -11316}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011100; Y = 8'b10000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 431,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11316
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000100; Y = 8'b00000111; // Expected: {'Z': -420}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000100; Y = 8'b00000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 432,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100110; Y = 8'b01101111; // Expected: {'Z': 4218}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100110; Y = 8'b01101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 433,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100011; Y = 8'b10101010; // Expected: {'Z': -3010}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100011; Y = 8'b10101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 434,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3010
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b10001010; // Expected: {'Z': -14514}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b10001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 435,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -14514
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110010; Y = 8'b11110001; // Expected: {'Z': -1710}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110010; Y = 8'b11110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 436,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1710
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b01110000; // Expected: {'Z': 4368}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b01110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 437,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000001; Y = 8'b11101100; // Expected: {'Z': -20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000001; Y = 8'b11101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 438,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010111; Y = 8'b00101111; // Expected: {'Z': 1081}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010111; Y = 8'b00101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 439,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1081
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b00001010; // Expected: {'Z': 680}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b00001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 440,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001000; Y = 8'b11101110; // Expected: {'Z': 2160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001000; Y = 8'b11101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 441,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b10111111; // Expected: {'Z': -4810}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b10111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 442,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4810
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100101; Y = 8'b10111010; // Expected: {'Z': 6370}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100101; Y = 8'b10111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 443,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6370
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b01011000; // Expected: {'Z': 4136}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b01011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 444,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011111; Y = 8'b11100011; // Expected: {'Z': -899}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011111; Y = 8'b11100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 445,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -899
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110000; Y = 8'b01100001; // Expected: {'Z': -7760}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110000; Y = 8'b01100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 446,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111000; Y = 8'b11100011; // Expected: {'Z': 2088}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111000; Y = 8'b11100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 447,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2088
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b11001111; // Expected: {'Z': -4704}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b11001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 448,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4704
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010001; Y = 8'b10010100; // Expected: {'Z': 5076}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010001; Y = 8'b10010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 449,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5076
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010010; Y = 8'b11101101; // Expected: {'Z': -342}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010010; Y = 8'b11101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 450,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -342
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111010; Y = 8'b01111111; // Expected: {'Z': 15494}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111010; Y = 8'b01111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 451,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 15494
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111111; Y = 8'b10011010; // Expected: {'Z': -6426}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111111; Y = 8'b10011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 452,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6426
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010100; Y = 8'b10010110; // Expected: {'Z': -8904}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010100; Y = 8'b10010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 453,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8904
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000001; Y = 8'b11001110; // Expected: {'Z': -3250}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000001; Y = 8'b11001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 454,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011101; Y = 8'b00110110; // Expected: {'Z': -5346}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011101; Y = 8'b00110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 455,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5346
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b11010000; // Expected: {'Z': -1008}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b11010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 456,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100011; Y = 8'b10000110; // Expected: {'Z': -4270}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100011; Y = 8'b10000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 457,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4270
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110001; Y = 8'b11111111; // Expected: {'Z': -113}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110001; Y = 8'b11111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 458,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110011; Y = 8'b00100101; // Expected: {'Z': 4255}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110011; Y = 8'b00100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 459,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011111; Y = 8'b01001111; // Expected: {'Z': -7663}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011111; Y = 8'b01001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 460,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7663
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b11111001; // Expected: {'Z': 609}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b11111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 461,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 609
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100111; Y = 8'b11001000; // Expected: {'Z': 1400}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100111; Y = 8'b11001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 462,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001010; Y = 8'b00011000; // Expected: {'Z': -2832}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001010; Y = 8'b00011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 463,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2832
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111011; Y = 8'b10100101; // Expected: {'Z': 6279}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111011; Y = 8'b10100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 464,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6279
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b11101101; // Expected: {'Z': 532}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b11101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 465,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 532
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011111; Y = 8'b01100011; // Expected: {'Z': 3069}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011111; Y = 8'b01100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 466,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3069
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011101; Y = 8'b00000001; // Expected: {'Z': -35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011101; Y = 8'b00000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 467,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010010; Y = 8'b11100100; // Expected: {'Z': 3080}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010010; Y = 8'b11100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 468,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010101; Y = 8'b00000110; // Expected: {'Z': -258}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010101; Y = 8'b00000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 469,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -258
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b01001011; // Expected: {'Z': -4425}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b01001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 470,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4425
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011000; Y = 8'b01111111; // Expected: {'Z': -5080}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011000; Y = 8'b01111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 471,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010111; Y = 8'b10011000; // Expected: {'Z': 10920}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010111; Y = 8'b10011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 472,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011001; Y = 8'b10000101; // Expected: {'Z': -10947}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011001; Y = 8'b10000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 473,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10947
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110101; Y = 8'b00100110; // Expected: {'Z': 4446}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110101; Y = 8'b00100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 474,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4446
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001111; Y = 8'b00010101; // Expected: {'Z': -2373}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001111; Y = 8'b00010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 475,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2373
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111010; Y = 8'b10110011; // Expected: {'Z': -4466}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111010; Y = 8'b10110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 476,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4466
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100011; Y = 8'b11100000; // Expected: {'Z': -1120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100011; Y = 8'b11100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 477,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100110; Y = 8'b11101100; // Expected: {'Z': 520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100110; Y = 8'b11101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 478,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011110; Y = 8'b11011011; // Expected: {'Z': -1110}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011110; Y = 8'b11011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 479,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011000; Y = 8'b01010000; // Expected: {'Z': 1920}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011000; Y = 8'b01010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 480,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101111; Y = 8'b11101000; // Expected: {'Z': 1944}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101111; Y = 8'b11101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 481,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111010; Y = 8'b10000000; // Expected: {'Z': 8960}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111010; Y = 8'b10000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 482,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100001; Y = 8'b11100001; // Expected: {'Z': 2945}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100001; Y = 8'b11100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 483,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2945
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001101; Y = 8'b01010110; // Expected: {'Z': 6622}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001101; Y = 8'b01010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 484,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6622
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b01001000; // Expected: {'Z': 648}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b01001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 485,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101000; Y = 8'b11010111; // Expected: {'Z': -1640}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101000; Y = 8'b11010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 486,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010000; Y = 8'b10010010; // Expected: {'Z': -8800}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010000; Y = 8'b10010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 487,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011111; Y = 8'b00101011; // Expected: {'Z': 1333}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011111; Y = 8'b00101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 488,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1333
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000011; Y = 8'b01011011; // Expected: {'Z': -5551}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000011; Y = 8'b01011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 489,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5551
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011010; Y = 8'b01100010; // Expected: {'Z': -9996}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011010; Y = 8'b01100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 490,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9996
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111100; Y = 8'b11011010; // Expected: {'Z': 152}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111100; Y = 8'b11011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 491,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100011; Y = 8'b01010101; // Expected: {'Z': -2465}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100011; Y = 8'b01010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 492,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2465
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b01111010; // Expected: {'Z': 2684}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b01111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 493,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2684
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100010; Y = 8'b01010011; // Expected: {'Z': 2822}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100010; Y = 8'b01010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 494,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2822
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101011; Y = 8'b00011011; // Expected: {'Z': 2889}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101011; Y = 8'b00011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 495,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2889
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101100; Y = 8'b00111110; // Expected: {'Z': 6696}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101100; Y = 8'b00111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 496,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6696
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011100; Y = 8'b00001000; // Expected: {'Z': 736}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011100; Y = 8'b00001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 497,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b10111000; // Expected: {'Z': -4392}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b10111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 498,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110100; Y = 8'b00100110; // Expected: {'Z': 4408}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110100; Y = 8'b00100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 499,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b00011010; // Expected: {'Z': -1456}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b00011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 500,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110010; Y = 8'b11001101; // Expected: {'Z': 714}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110010; Y = 8'b11001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 501,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 714
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100011; Y = 8'b10010011; // Expected: {'Z': 3161}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100011; Y = 8'b10010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 502,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3161
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010010; Y = 8'b11011111; // Expected: {'Z': -594}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010010; Y = 8'b11011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 503,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -594
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000101; Y = 8'b11000100; // Expected: {'Z': 7380}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000101; Y = 8'b11000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 504,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7380
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110100; Y = 8'b11101100; // Expected: {'Z': -1040}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110100; Y = 8'b11101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 505,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001110; Y = 8'b11101110; // Expected: {'Z': 2052}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001110; Y = 8'b11101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 506,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2052
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110010; Y = 8'b01011001; // Expected: {'Z': 10146}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110010; Y = 8'b01011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 507,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000011; Y = 8'b10010100; // Expected: {'Z': 6588}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000011; Y = 8'b10010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 508,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6588
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101001; Y = 8'b10100001; // Expected: {'Z': -3895}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101001; Y = 8'b10100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 509,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3895
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101111; Y = 8'b10101010; // Expected: {'Z': -9546}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101111; Y = 8'b10101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 510,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011110; Y = 8'b11111011; // Expected: {'Z': 170}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011110; Y = 8'b11111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 511,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101010; Y = 8'b01011110; // Expected: {'Z': -8084}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101010; Y = 8'b01011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 512,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8084
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100110; Y = 8'b00100010; // Expected: {'Z': 3468}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100110; Y = 8'b00100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 513,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3468
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100000; Y = 8'b10001110; // Expected: {'Z': 3648}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100000; Y = 8'b10001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 514,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010011; Y = 8'b10000101; // Expected: {'Z': 5535}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010011; Y = 8'b10000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 515,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5535
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111010; Y = 8'b00110110; // Expected: {'Z': 6588}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111010; Y = 8'b00110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 516,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6588
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000111; Y = 8'b10010010; // Expected: {'Z': -7810}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000111; Y = 8'b10010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 517,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7810
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111011; Y = 8'b11010110; // Expected: {'Z': -2478}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111011; Y = 8'b11010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 518,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2478
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b01111101; // Expected: {'Z': 12000}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b01111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 519,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 12000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110010; Y = 8'b10110010; // Expected: {'Z': -3900}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110010; Y = 8'b10110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 520,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001001; Y = 8'b01110010; // Expected: {'Z': -13566}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001001; Y = 8'b01110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 521,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -13566
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111010; Y = 8'b10001001; // Expected: {'Z': -6902}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111010; Y = 8'b10001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 522,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6902
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100101; Y = 8'b10101000; // Expected: {'Z': 2376}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100101; Y = 8'b10101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 523,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2376
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101001; Y = 8'b00101110; // Expected: {'Z': -1058}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101001; Y = 8'b00101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 524,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1058
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000101; Y = 8'b11010110; // Expected: {'Z': -210}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000101; Y = 8'b11010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 525,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b11110011; // Expected: {'Z': -78}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b11110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 526,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001110; Y = 8'b10001100; // Expected: {'Z': -1624}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001110; Y = 8'b10001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 527,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010010; Y = 8'b11100001; // Expected: {'Z': 1426}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010010; Y = 8'b11100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 528,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1426
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b11000111; // Expected: {'Z': -3477}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b11000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 529,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3477
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010011; Y = 8'b01011000; // Expected: {'Z': 7304}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010011; Y = 8'b01011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 530,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7304
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100011; Y = 8'b00010111; // Expected: {'Z': -667}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100011; Y = 8'b00010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 531,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -667
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001101; Y = 8'b11111111; // Expected: {'Z': 115}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001101; Y = 8'b11111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 532,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 115
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100011; Y = 8'b01001011; // Expected: {'Z': -2175}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100011; Y = 8'b01001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 533,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000011; Y = 8'b01111110; // Expected: {'Z': 378}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000011; Y = 8'b01111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 534,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 378
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010010; Y = 8'b00011111; // Expected: {'Z': 558}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010010; Y = 8'b00011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 535,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 558
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011000; Y = 8'b10000010; // Expected: {'Z': -3024}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011000; Y = 8'b10000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 536,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100000; Y = 8'b01010000; // Expected: {'Z': 2560}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100000; Y = 8'b01010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 537,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010011; Y = 8'b00110100; // Expected: {'Z': 4316}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010011; Y = 8'b00110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 538,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4316
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b11100101; // Expected: {'Z': 2997}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b11100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 539,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2997
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111100; Y = 8'b10001001; // Expected: {'Z': 476}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111100; Y = 8'b10001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 540,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 476
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111101; Y = 8'b11110011; // Expected: {'Z': -1625}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111101; Y = 8'b11110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 541,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1625
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011100; Y = 8'b11100000; // Expected: {'Z': 1152}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011100; Y = 8'b11100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 542,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b10100011; // Expected: {'Z': 5208}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b10100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 543,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100011; Y = 8'b00110110; // Expected: {'Z': 1890}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100011; Y = 8'b00110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 544,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1890
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010000; Y = 8'b10010111; // Expected: {'Z': 5040}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010000; Y = 8'b10010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 545,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b11100110; // Expected: {'Z': -2496}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b11100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 546,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110011; Y = 8'b00101111; // Expected: {'Z': -3619}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110011; Y = 8'b00101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 547,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3619
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b11110100; // Expected: {'Z': -108}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b11110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 548,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110100; Y = 8'b10100001; // Expected: {'Z': -11020}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110100; Y = 8'b10100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 549,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11020
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100011; Y = 8'b10011101; // Expected: {'Z': 2871}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100011; Y = 8'b10011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 550,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2871
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010101; Y = 8'b00100100; // Expected: {'Z': -3852}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010101; Y = 8'b00100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 551,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3852
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001100; Y = 8'b00000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001100; Y = 8'b00000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 552,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111111; Y = 8'b01001001; // Expected: {'Z': -73}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111111; Y = 8'b01001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 553,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110110; Y = 8'b11111110; // Expected: {'Z': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110110; Y = 8'b11111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 554,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b10011111; // Expected: {'Z': -2037}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b10011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 555,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2037
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011110; Y = 8'b01110111; // Expected: {'Z': 3570}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011110; Y = 8'b01110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 556,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3570
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101001; Y = 8'b00010000; // Expected: {'Z': -368}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101001; Y = 8'b00010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 557,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100000; Y = 8'b11110010; // Expected: {'Z': 448}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100000; Y = 8'b11110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 558,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 448
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011001; Y = 8'b00001000; // Expected: {'Z': -824}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011001; Y = 8'b00001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 559,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -824
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101011; Y = 8'b11100101; // Expected: {'Z': 567}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101011; Y = 8'b11100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 560,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 567
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001110; Y = 8'b00011101; // Expected: {'Z': -3306}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001110; Y = 8'b00011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 561,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3306
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001010; Y = 8'b11011010; // Expected: {'Z': 4484}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001010; Y = 8'b11011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 562,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4484
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b01111000; // Expected: {'Z': 2640}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b01111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 563,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100011; Y = 8'b00101110; // Expected: {'Z': 4554}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100011; Y = 8'b00101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 564,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4554
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011011; Y = 8'b11101011; // Expected: {'Z': 2121}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011011; Y = 8'b11101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 565,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011000; Y = 8'b01010101; // Expected: {'Z': -3400}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011000; Y = 8'b01010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 566,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b11010110; // Expected: {'Z': 3528}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b11010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 567,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111001; Y = 8'b10101110; // Expected: {'Z': 5822}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111001; Y = 8'b10101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 568,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5822
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b11000000; // Expected: {'Z': -1344}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b11000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 569,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1344
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110011; Y = 8'b01000110; // Expected: {'Z': 8050}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110011; Y = 8'b01000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 570,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011101; Y = 8'b11110000; // Expected: {'Z': -1488}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011101; Y = 8'b11110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 571,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111011; Y = 8'b11111111; // Expected: {'Z': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111011; Y = 8'b11111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 572,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b10110110; // Expected: {'Z': -7104}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b10110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 573,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111011; Y = 8'b11110011; // Expected: {'Z': 65}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111011; Y = 8'b11110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 574,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b00011100; // Expected: {'Z': 1708}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b00011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 575,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1708
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110110; Y = 8'b10010111; // Expected: {'Z': -12390}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110110; Y = 8'b10010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 576,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12390
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110111; Y = 8'b10101001; // Expected: {'Z': 783}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110111; Y = 8'b10101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 577,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 783
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111000; Y = 8'b11110001; // Expected: {'Z': -1800}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111000; Y = 8'b11110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 578,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000101; Y = 8'b11110100; // Expected: {'Z': 1476}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000101; Y = 8'b11110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 579,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1476
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110111; Y = 8'b11111111; // Expected: {'Z': -55}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110111; Y = 8'b11111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 580,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b00010100; // Expected: {'Z': 260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b00010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 581,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b01001111; // Expected: {'Z': 1185}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b01001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 582,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010111; Y = 8'b01110101; // Expected: {'Z': 10179}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010111; Y = 8'b01110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 583,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10179
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011110; Y = 8'b11100010; // Expected: {'Z': -2820}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011110; Y = 8'b11100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 584,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b01010101; // Expected: {'Z': 6290}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b01010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 585,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6290
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001010; Y = 8'b00010001; // Expected: {'Z': -2006}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001010; Y = 8'b00010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 586,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2006
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011010; Y = 8'b10100001; // Expected: {'Z': -2470}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011010; Y = 8'b10100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 587,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2470
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010101; Y = 8'b10010100; // Expected: {'Z': -9180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010101; Y = 8'b10010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 588,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000001; Y = 8'b11000111; // Expected: {'Z': -3705}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000001; Y = 8'b11000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 589,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3705
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101101; Y = 8'b11000000; // Expected: {'Z': -2880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101101; Y = 8'b11000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 590,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010001; Y = 8'b10110110; // Expected: {'Z': -5994}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010001; Y = 8'b10110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 591,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5994
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b10100011; // Expected: {'Z': 10323}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b10100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 592,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10323
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b11100000; // Expected: {'Z': 2784}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b11100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 593,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011100; Y = 8'b10010100; // Expected: {'Z': 3888}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011100; Y = 8'b10010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 594,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110111; Y = 8'b10010011; // Expected: {'Z': 7957}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110111; Y = 8'b10010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 595,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7957
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010111; Y = 8'b11101111; // Expected: {'Z': 1785}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010111; Y = 8'b11101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 596,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1785
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101110; Y = 8'b00100110; // Expected: {'Z': 4180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101110; Y = 8'b00100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 597,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010111; Y = 8'b01010000; // Expected: {'Z': 6960}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010111; Y = 8'b01010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 598,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111011; Y = 8'b11010001; // Expected: {'Z': -2773}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111011; Y = 8'b11010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 599,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2773
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110110; Y = 8'b01000000; // Expected: {'Z': -640}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110110; Y = 8'b01000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 600,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011101; Y = 8'b00000001; // Expected: {'Z': 93}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011101; Y = 8'b00000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 601,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000100; Y = 8'b01110000; // Expected: {'Z': -13888}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000100; Y = 8'b01110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 602,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -13888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000100; Y = 8'b01110010; // Expected: {'Z': -6840}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000100; Y = 8'b01110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 603,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100011; Y = 8'b01001011; // Expected: {'Z': -2175}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100011; Y = 8'b01001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 604,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101011; Y = 8'b10001000; // Expected: {'Z': -5160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101011; Y = 8'b10001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 605,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b10100110; // Expected: {'Z': -1710}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b10100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 606,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1710
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011001; Y = 8'b00010101; // Expected: {'Z': 1869}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011001; Y = 8'b00010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 607,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1869
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b10001111; // Expected: {'Z': -2373}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b10001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 608,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2373
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b01101001; // Expected: {'Z': 945}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b01101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 609,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 945
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b01001010; // Expected: {'Z': 1110}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b01001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 610,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010101; Y = 8'b11100101; // Expected: {'Z': 1161}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010101; Y = 8'b11100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 611,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1161
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001100; Y = 8'b11101010; // Expected: {'Z': -264}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001100; Y = 8'b11101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 612,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111001; Y = 8'b01011010; // Expected: {'Z': -6390}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111001; Y = 8'b01011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 613,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6390
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101010; Y = 8'b10011010; // Expected: {'Z': 8772}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101010; Y = 8'b10011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 614,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8772
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111010; Y = 8'b00010101; // Expected: {'Z': 1218}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111010; Y = 8'b00010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 615,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b10100000; // Expected: {'Z': 8352}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b10100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 616,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b11000110; // Expected: {'Z': -754}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b11000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 617,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -754
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000011; Y = 8'b10001111; // Expected: {'Z': -7571}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000011; Y = 8'b10001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 618,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7571
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100110; Y = 8'b00010100; // Expected: {'Z': -520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100110; Y = 8'b00010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 619,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111000; Y = 8'b10111110; // Expected: {'Z': 4752}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111000; Y = 8'b10111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 620,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4752
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110101; Y = 8'b00100010; // Expected: {'Z': -2550}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110101; Y = 8'b00100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 621,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000000; Y = 8'b11110111; // Expected: {'Z': 576}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000000; Y = 8'b11110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 622,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000011; Y = 8'b10000011; // Expected: {'Z': 15625}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000011; Y = 8'b10000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 623,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 15625
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000100; Y = 8'b00111110; // Expected: {'Z': -7688}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000100; Y = 8'b00111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 624,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7688
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b01101111; // Expected: {'Z': 11433}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b01101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 625,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11433
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011100; Y = 8'b01100001; // Expected: {'Z': -3492}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011100; Y = 8'b01100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 626,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3492
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000111; Y = 8'b11000011; // Expected: {'Z': -427}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000111; Y = 8'b11000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 627,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -427
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111110; Y = 8'b11010100; // Expected: {'Z': 2904}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111110; Y = 8'b11010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 628,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2904
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001110; Y = 8'b00100000; // Expected: {'Z': -1600}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001110; Y = 8'b00100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 629,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001110; Y = 8'b01111110; // Expected: {'Z': -6300}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001110; Y = 8'b01111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 630,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100000; Y = 8'b00010001; // Expected: {'Z': -1632}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100000; Y = 8'b00010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 631,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1632
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010111; Y = 8'b10001010; // Expected: {'Z': -2714}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010111; Y = 8'b10001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 632,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2714
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101010; Y = 8'b01110100; // Expected: {'Z': 12296}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101010; Y = 8'b01110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 633,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 12296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010100; Y = 8'b10110001; // Expected: {'Z': -1580}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010100; Y = 8'b10110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 634,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100110; Y = 8'b01101010; // Expected: {'Z': -2756}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100110; Y = 8'b01101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 635,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b00000100; // Expected: {'Z': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b00000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 636,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100101; Y = 8'b10110100; // Expected: {'Z': -2812}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100101; Y = 8'b10110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 637,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2812
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b11000111; // Expected: {'Z': -4218}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b11000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 638,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011010; Y = 8'b10001000; // Expected: {'Z': 12240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011010; Y = 8'b10001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 639,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 12240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b00101100; // Expected: {'Z': 836}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b00101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 640,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 836
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b11010001; // Expected: {'Z': 2632}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b11010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 641,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2632
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b01000100; // Expected: {'Z': 1496}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b01000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 642,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100100; Y = 8'b11110101; // Expected: {'Z': 1012}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100100; Y = 8'b11110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 643,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1012
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101011; Y = 8'b00110000; // Expected: {'Z': -4080}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101011; Y = 8'b00110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 644,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111111; Y = 8'b00011101; // Expected: {'Z': -1885}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111111; Y = 8'b00011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 645,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1885
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101001; Y = 8'b10010011; // Expected: {'Z': 2507}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101001; Y = 8'b10010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 646,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2507
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111100; Y = 8'b10111001; // Expected: {'Z': -4260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111100; Y = 8'b10111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 647,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010001; Y = 8'b11010010; // Expected: {'Z': -3726}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010001; Y = 8'b11010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 648,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3726
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000111; Y = 8'b11001011; // Expected: {'Z': 3021}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000111; Y = 8'b11001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 649,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3021
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101101; Y = 8'b11100111; // Expected: {'Z': 475}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101101; Y = 8'b11100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 650,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 475
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011111; Y = 8'b00001110; // Expected: {'Z': 1330}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011111; Y = 8'b00001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 651,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1330
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111100; Y = 8'b10100111; // Expected: {'Z': -5340}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111100; Y = 8'b10100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 652,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000000; Y = 8'b00100111; // Expected: {'Z': -4992}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000000; Y = 8'b00100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 653,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4992
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001110; Y = 8'b11010110; // Expected: {'Z': 4788}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001110; Y = 8'b11010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 654,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4788
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101001; Y = 8'b00111111; // Expected: {'Z': 6615}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101001; Y = 8'b00111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 655,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6615
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011001; Y = 8'b10101100; // Expected: {'Z': -2100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011001; Y = 8'b10101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 656,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b00111011; // Expected: {'Z': 2773}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b00111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 657,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2773
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001000; Y = 8'b01000111; // Expected: {'Z': -8520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001000; Y = 8'b01000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 658,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010010; Y = 8'b01111100; // Expected: {'Z': -13640}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010010; Y = 8'b01111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 659,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -13640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b00001111; // Expected: {'Z': 1110}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b00001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 660,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011010; Y = 8'b01010010; // Expected: {'Z': -3116}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011010; Y = 8'b01010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 661,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b01101110; // Expected: {'Z': 2090}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b01101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 662,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2090
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010001; Y = 8'b00001010; // Expected: {'Z': -470}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010001; Y = 8'b00001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 663,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -470
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000011; Y = 8'b01001000; // Expected: {'Z': 4824}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000011; Y = 8'b01001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 664,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4824
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001110; Y = 8'b11110000; // Expected: {'Z': 800}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001110; Y = 8'b11110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 665,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101100; Y = 8'b11010101; // Expected: {'Z': -4644}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101100; Y = 8'b11010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 666,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4644
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b10101101; // Expected: {'Z': -498}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b10101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 667,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -498
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100100; Y = 8'b01110000; // Expected: {'Z': 11200}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100100; Y = 8'b01110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 668,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101101; Y = 8'b10101111; // Expected: {'Z': 6723}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101101; Y = 8'b10101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 669,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6723
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b11011001; // Expected: {'Z': -1131}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b11011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 670,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111100; Y = 8'b11010010; // Expected: {'Z': -2760}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111100; Y = 8'b11010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 671,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010100; Y = 8'b10110010; // Expected: {'Z': -6552}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010100; Y = 8'b10110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 672,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010110; Y = 8'b10000011; // Expected: {'Z': 13250}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010110; Y = 8'b10000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 673,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 13250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011100; Y = 8'b00010011; // Expected: {'Z': -1900}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011100; Y = 8'b00010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 674,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110011; Y = 8'b11001101; // Expected: {'Z': -5865}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110011; Y = 8'b11001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 675,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5865
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101111; Y = 8'b10110000; // Expected: {'Z': 6480}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101111; Y = 8'b10110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 676,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101010; Y = 8'b10100101; // Expected: {'Z': -3822}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101010; Y = 8'b10100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 677,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3822
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111100; Y = 8'b10001000; // Expected: {'Z': -7200}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111100; Y = 8'b10001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 678,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110101; Y = 8'b11100110; // Expected: {'Z': -3042}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110101; Y = 8'b11100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 679,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3042
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110000; Y = 8'b10100101; // Expected: {'Z': -4368}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110000; Y = 8'b10100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 680,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100110; Y = 8'b10110011; // Expected: {'Z': -7854}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100110; Y = 8'b10110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 681,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7854
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100100; Y = 8'b00100100; // Expected: {'Z': 3600}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100100; Y = 8'b00100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 682,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011111; Y = 8'b01100001; // Expected: {'Z': -9409}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011111; Y = 8'b01100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 683,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9409
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b00100000; // Expected: {'Z': -2176}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b00100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 684,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b10010110; // Expected: {'Z': -2226}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b10010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 685,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2226
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111011; Y = 8'b10001101; // Expected: {'Z': 7935}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111011; Y = 8'b10001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 686,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7935
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000011; Y = 8'b10111110; // Expected: {'Z': -4422}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000011; Y = 8'b10111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 687,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4422
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110000; Y = 8'b00001010; // Expected: {'Z': -800}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110000; Y = 8'b00001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 688,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000000; Y = 8'b00001100; // Expected: {'Z': -1536}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000000; Y = 8'b00001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 689,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1536
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000111; Y = 8'b00011000; // Expected: {'Z': -1368}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000111; Y = 8'b00011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 690,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011011; Y = 8'b01101011; // Expected: {'Z': -10807}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011011; Y = 8'b01101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 691,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10807
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011110; Y = 8'b00000001; // Expected: {'Z': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011110; Y = 8'b00000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 692,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b00001110; // Expected: {'Z': -784}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b00001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 693,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100111; Y = 8'b10011011; // Expected: {'Z': 8989}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100111; Y = 8'b10011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 694,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8989
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111110; Y = 8'b00111101; // Expected: {'Z': -122}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111110; Y = 8'b00111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 695,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101010; Y = 8'b10111001; // Expected: {'Z': -7526}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101010; Y = 8'b10111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 696,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7526
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011111; Y = 8'b11100001; // Expected: {'Z': 3007}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011111; Y = 8'b11100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 697,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3007
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110101; Y = 8'b01010010; // Expected: {'Z': 9594}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110101; Y = 8'b01010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 698,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9594
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011101; Y = 8'b00001011; // Expected: {'Z': -385}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011101; Y = 8'b00001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 699,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -385
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110110; Y = 8'b11010011; // Expected: {'Z': 450}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110110; Y = 8'b11010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 700,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b00001110; // Expected: {'Z': 1232}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b00001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 701,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101001; Y = 8'b00001011; // Expected: {'Z': 451}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101001; Y = 8'b00001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 702,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 451
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100001; Y = 8'b11100101; // Expected: {'Z': -2619}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100001; Y = 8'b11100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 703,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2619
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b00001011; // Expected: {'Z': 594}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b00001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 704,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 594
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111111; Y = 8'b10110011; // Expected: {'Z': -4851}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111111; Y = 8'b10110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 705,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4851
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101111; Y = 8'b10101001; // Expected: {'Z': 7047}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101111; Y = 8'b10101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 706,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7047
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111010; Y = 8'b01010100; // Expected: {'Z': 10248}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111010; Y = 8'b01010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 707,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110000; Y = 8'b11001101; // Expected: {'Z': 816}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110000; Y = 8'b11001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 708,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100111; Y = 8'b11000110; // Expected: {'Z': 1450}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100111; Y = 8'b11000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 709,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111001; Y = 8'b10001010; // Expected: {'Z': 8378}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111001; Y = 8'b10001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 710,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8378
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001001; Y = 8'b11100010; // Expected: {'Z': -2190}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001001; Y = 8'b11100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 711,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110101; Y = 8'b10101011; // Expected: {'Z': -9945}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110101; Y = 8'b10101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 712,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9945
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111000; Y = 8'b01100000; // Expected: {'Z': -768}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111000; Y = 8'b01100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 713,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -768
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010001; Y = 8'b01101000; // Expected: {'Z': 1768}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010001; Y = 8'b01101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 714,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1768
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b01101000; // Expected: {'Z': -9048}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b01101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 715,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9048
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b10110000; // Expected: {'Z': 6960}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b10110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 716,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b11010010; // Expected: {'Z': -3312}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b11010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 717,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3312
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011011; Y = 8'b10101000; // Expected: {'Z': 3256}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011011; Y = 8'b10101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 718,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3256
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110010; Y = 8'b10001010; // Expected: {'Z': -13452}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110010; Y = 8'b10001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 719,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -13452
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111000; Y = 8'b01011001; // Expected: {'Z': -712}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111000; Y = 8'b01011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 720,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -712
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101000; Y = 8'b10001101; // Expected: {'Z': -4600}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101000; Y = 8'b10001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 721,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010110; Y = 8'b11001110; // Expected: {'Z': 5300}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010110; Y = 8'b11001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 722,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001010; Y = 8'b11001111; // Expected: {'Z': -490}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001010; Y = 8'b11001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 723,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -490
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001011; Y = 8'b00010000; // Expected: {'Z': 1200}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001011; Y = 8'b00010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 724,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000000; Y = 8'b01011010; // Expected: {'Z': -11520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000000; Y = 8'b01011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 725,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100001; Y = 8'b10111000; // Expected: {'Z': 2232}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100001; Y = 8'b10111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 726,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111001; Y = 8'b11111011; // Expected: {'Z': 355}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111001; Y = 8'b11111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 727,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 355
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b10100110; // Expected: {'Z': 4590}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b10100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 728,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4590
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b01101110; // Expected: {'Z': 13530}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b01101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 729,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 13530
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111101; Y = 8'b10000000; // Expected: {'Z': -16000}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111101; Y = 8'b10000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 730,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -16000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110010; Y = 8'b01000101; // Expected: {'Z': 7866}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110010; Y = 8'b01000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 731,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7866
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110011; Y = 8'b11000000; // Expected: {'Z': 832}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110011; Y = 8'b11000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 732,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 832
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010000; Y = 8'b00110010; // Expected: {'Z': 4000}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010000; Y = 8'b00110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 733,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110111; Y = 8'b11000010; // Expected: {'Z': -7378}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110111; Y = 8'b11000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 734,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7378
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100101; Y = 8'b10000101; // Expected: {'Z': 3321}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100101; Y = 8'b10000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 735,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3321
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000010; Y = 8'b11101000; // Expected: {'Z': -1584}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000010; Y = 8'b11101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 736,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1584
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110111; Y = 8'b10000010; // Expected: {'Z': 1134}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110111; Y = 8'b10000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 737,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110111; Y = 8'b11000100; // Expected: {'Z': -3300}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110111; Y = 8'b11000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 738,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101010; Y = 8'b01101101; // Expected: {'Z': 4578}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101010; Y = 8'b01101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 739,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4578
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101111; Y = 8'b11110110; // Expected: {'Z': -1110}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101111; Y = 8'b11110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 740,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b01111000; // Expected: {'Z': -7080}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b01111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 741,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000010; Y = 8'b01001111; // Expected: {'Z': 5214}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000010; Y = 8'b01001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 742,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111000; Y = 8'b10111010; // Expected: {'Z': 560}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111000; Y = 8'b10111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 743,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001001; Y = 8'b10001100; // Expected: {'Z': -8468}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001001; Y = 8'b10001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 744,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8468
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010101; Y = 8'b01101100; // Expected: {'Z': -4644}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010101; Y = 8'b01101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 745,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4644
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000000; Y = 8'b11110101; // Expected: {'Z': 1408}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000000; Y = 8'b11110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 746,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101100; Y = 8'b01010010; // Expected: {'Z': -1640}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101100; Y = 8'b01010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 747,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010111; Y = 8'b10011000; // Expected: {'Z': -9048}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010111; Y = 8'b10011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 748,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9048
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b11000011; // Expected: {'Z': 6771}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b11000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 749,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6771
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101011; Y = 8'b01000000; // Expected: {'Z': 6848}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101011; Y = 8'b01000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 750,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b10001101; // Expected: {'Z': -11845}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b10001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 751,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11845
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010111; Y = 8'b10001110; // Expected: {'Z': 4674}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010111; Y = 8'b10001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 752,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4674
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010010; Y = 8'b01000000; // Expected: {'Z': 1152}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010010; Y = 8'b01000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 753,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010100; Y = 8'b01011110; // Expected: {'Z': -4136}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010100; Y = 8'b01011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 754,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001011; Y = 8'b00011111; // Expected: {'Z': -1643}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001011; Y = 8'b00011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 755,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1643
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011001; Y = 8'b10101101; // Expected: {'Z': 3237}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011001; Y = 8'b10101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 756,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3237
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101101; Y = 8'b00110110; // Expected: {'Z': 2430}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101101; Y = 8'b00110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 757,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110010; Y = 8'b11111011; // Expected: {'Z': 70}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110010; Y = 8'b11111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 758,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001000; Y = 8'b01000110; // Expected: {'Z': -8400}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001000; Y = 8'b01000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 759,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100010; Y = 8'b00100100; // Expected: {'Z': 1224}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100010; Y = 8'b00100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 760,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010101; Y = 8'b11100011; // Expected: {'Z': 3103}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010101; Y = 8'b11100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 761,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b01111101; // Expected: {'Z': 3625}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b01111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 762,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3625
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001100; Y = 8'b10110101; // Expected: {'Z': -5700}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001100; Y = 8'b10110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 763,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101001; Y = 8'b11011110; // Expected: {'Z': -1394}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101001; Y = 8'b11011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 764,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1394
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010000; Y = 8'b01111100; // Expected: {'Z': -5952}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010000; Y = 8'b01111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 765,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5952
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111101; Y = 8'b11111001; // Expected: {'Z': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111101; Y = 8'b11111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 766,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000111; Y = 8'b11011110; // Expected: {'Z': 4114}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000111; Y = 8'b11011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 767,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b01011001; // Expected: {'Z': 3916}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b01011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 768,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3916
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001000; Y = 8'b10110100; // Expected: {'Z': 9120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001000; Y = 8'b10110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 769,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100101; Y = 8'b11111111; // Expected: {'Z': -101}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100101; Y = 8'b11111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 770,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011001; Y = 8'b10010011; // Expected: {'Z': -2725}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011001; Y = 8'b10010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 771,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2725
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101100; Y = 8'b11100011; // Expected: {'Z': -3132}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101100; Y = 8'b11100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 772,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100110; Y = 8'b11110001; // Expected: {'Z': 1350}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100110; Y = 8'b11110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 773,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001111; Y = 8'b01010110; // Expected: {'Z': -9718}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001111; Y = 8'b01010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 774,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9718
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001000; Y = 8'b11001111; // Expected: {'Z': -392}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001000; Y = 8'b11001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 775,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b01001011; // Expected: {'Z': 9225}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b01001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 776,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111110; Y = 8'b10111111; // Expected: {'Z': -4030}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111110; Y = 8'b10111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 777,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4030
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b11111010; // Expected: {'Z': -216}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b11111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 778,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110100; Y = 8'b10111010; // Expected: {'Z': -8120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110100; Y = 8'b10111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 779,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010100; Y = 8'b01000100; // Expected: {'Z': 5712}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010100; Y = 8'b01000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 780,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5712
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001000; Y = 8'b00110000; // Expected: {'Z': 384}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001000; Y = 8'b00110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 781,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 384
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110110; Y = 8'b01000100; // Expected: {'Z': -680}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110110; Y = 8'b01000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 782,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111011; Y = 8'b10011000; // Expected: {'Z': 520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111011; Y = 8'b10011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 783,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b10111111; // Expected: {'Z': 5330}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b10111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 784,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5330
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010111; Y = 8'b00010101; // Expected: {'Z': 483}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010111; Y = 8'b00010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 785,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 483
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001110; Y = 8'b10100001; // Expected: {'Z': 10830}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001110; Y = 8'b10100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 786,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10830
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101001; Y = 8'b11111011; // Expected: {'Z': -525}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101001; Y = 8'b11111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 787,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -525
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000111; Y = 8'b01101110; // Expected: {'Z': 7810}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000111; Y = 8'b01101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 788,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7810
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001111; Y = 8'b00011101; // Expected: {'Z': -3277}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001111; Y = 8'b00011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 789,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3277
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100100; Y = 8'b01100000; // Expected: {'Z': -8832}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100100; Y = 8'b01100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 790,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8832
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001001; Y = 8'b00011111; // Expected: {'Z': -1705}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001001; Y = 8'b00011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 791,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1705
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001110; Y = 8'b01000001; // Expected: {'Z': 910}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001110; Y = 8'b01000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 792,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 910
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b01010010; // Expected: {'Z': 3198}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b01010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 793,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011101; Y = 8'b00001000; // Expected: {'Z': 744}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011101; Y = 8'b00001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 794,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 744
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010110; Y = 8'b00101010; // Expected: {'Z': -4452}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010110; Y = 8'b00101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 795,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4452
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010110; Y = 8'b00101100; // Expected: {'Z': 3784}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010110; Y = 8'b00101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 796,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110001; Y = 8'b10011011; // Expected: {'Z': -4949}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110001; Y = 8'b10011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 797,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4949
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110010; Y = 8'b11000001; // Expected: {'Z': -7182}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110010; Y = 8'b11000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 798,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011000; Y = 8'b11001101; // Expected: {'Z': 2040}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011000; Y = 8'b11001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 799,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010111; Y = 8'b11101001; // Expected: {'Z': 2415}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010111; Y = 8'b11101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 800,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2415
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010010; Y = 8'b11101011; // Expected: {'Z': 2310}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010010; Y = 8'b11101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 801,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2310
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110111; Y = 8'b11010001; // Expected: {'Z': 3431}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110111; Y = 8'b11010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 802,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3431
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001110; Y = 8'b10011111; // Expected: {'Z': 11058}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001110; Y = 8'b10011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 803,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11058
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010001; Y = 8'b00111100; // Expected: {'Z': 4860}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010001; Y = 8'b00111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 804,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4860
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010100; Y = 8'b01100111; // Expected: {'Z': -11124}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010100; Y = 8'b01100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 805,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010100; Y = 8'b00011111; // Expected: {'Z': -3348}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010100; Y = 8'b00011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 806,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3348
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b11111000; // Expected: {'Z': -544}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b11111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 807,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -544
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111110; Y = 8'b00000111; // Expected: {'Z': -462}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111110; Y = 8'b00000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 808,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001101; Y = 8'b01101010; // Expected: {'Z': -12190}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001101; Y = 8'b01101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 809,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011101; Y = 8'b11110101; // Expected: {'Z': 385}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011101; Y = 8'b11110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 810,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 385
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110001; Y = 8'b00011001; // Expected: {'Z': 1225}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110001; Y = 8'b00011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 811,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001001; Y = 8'b10111110; // Expected: {'Z': 3630}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001001; Y = 8'b10111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 812,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3630
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011001; Y = 8'b00010000; // Expected: {'Z': 400}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011001; Y = 8'b00010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 813,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100010; Y = 8'b00011100; // Expected: {'Z': 952}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100010; Y = 8'b00011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 814,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 952
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011011; Y = 8'b01111011; // Expected: {'Z': -12423}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011011; Y = 8'b01111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 815,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12423
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110000; Y = 8'b00101111; // Expected: {'Z': 2256}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110000; Y = 8'b00101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 816,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2256
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001101; Y = 8'b11011101; // Expected: {'Z': 4025}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001101; Y = 8'b11011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 817,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4025
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000010; Y = 8'b01001011; // Expected: {'Z': 4950}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000010; Y = 8'b01001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 818,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011100; Y = 8'b10111101; // Expected: {'Z': -6164}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011100; Y = 8'b10111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 819,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000101; Y = 8'b11000011; // Expected: {'Z': -4209}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000101; Y = 8'b11000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 820,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010000; Y = 8'b10001000; // Expected: {'Z': 13440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010000; Y = 8'b10001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 821,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 13440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001000; Y = 8'b00001111; // Expected: {'Z': 120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001000; Y = 8'b00001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 822,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b10011110; // Expected: {'Z': -2842}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b10011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 823,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2842
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100000; Y = 8'b01101111; // Expected: {'Z': -3552}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100000; Y = 8'b01101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 824,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011101; Y = 8'b11010000; // Expected: {'Z': -4464}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011101; Y = 8'b11010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 825,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b11100100; // Expected: {'Z': -1316}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b11100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 826,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1316
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010100; Y = 8'b10100111; // Expected: {'Z': -7476}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010100; Y = 8'b10100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 827,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7476
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111011; Y = 8'b00000100; // Expected: {'Z': 236}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111011; Y = 8'b00000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 828,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001100; Y = 8'b11111100; // Expected: {'Z': -304}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001100; Y = 8'b11111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 829,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -304
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111010; Y = 8'b10010001; // Expected: {'Z': 7770}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111010; Y = 8'b10010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 830,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7770
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000100; Y = 8'b10011010; // Expected: {'Z': 6120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000100; Y = 8'b10011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 831,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b00111101; // Expected: {'Z': 6283}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b00111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 832,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6283
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010000; Y = 8'b00010010; // Expected: {'Z': -864}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010000; Y = 8'b00010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 833,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -864
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101000; Y = 8'b11010100; // Expected: {'Z': -1760}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101000; Y = 8'b11010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 834,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b01100000; // Expected: {'Z': -10656}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b01100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 835,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10656
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111010; Y = 8'b01000111; // Expected: {'Z': -426}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111010; Y = 8'b01000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 836,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -426
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111000; Y = 8'b01110010; // Expected: {'Z': 13680}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111000; Y = 8'b01110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 837,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 13680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b00010111; // Expected: {'Z': 506}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b00010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 838,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 506
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000011; Y = 8'b10000010; // Expected: {'Z': 7686}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000011; Y = 8'b10000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 839,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7686
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100011; Y = 8'b10001111; // Expected: {'Z': -3955}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100011; Y = 8'b10001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 840,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3955
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101011; Y = 8'b11001111; // Expected: {'Z': 1029}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101011; Y = 8'b11001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 841,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1029
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101011; Y = 8'b11000111; // Expected: {'Z': 4845}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101011; Y = 8'b11000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 842,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4845
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000110; Y = 8'b10111011; // Expected: {'Z': -4830}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000110; Y = 8'b10111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 843,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4830
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111011; Y = 8'b11110111; // Expected: {'Z': 45}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111011; Y = 8'b11110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 844,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b11000100; // Expected: {'Z': -5760}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b11000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 845,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101010; Y = 8'b10111011; // Expected: {'Z': 5934}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101010; Y = 8'b10111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 846,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5934
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100010; Y = 8'b11101101; // Expected: {'Z': -1862}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100010; Y = 8'b11101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 847,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1862
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110100; Y = 8'b10100100; // Expected: {'Z': 6992}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110100; Y = 8'b10100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 848,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6992
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010000; Y = 8'b00111110; // Expected: {'Z': 4960}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010000; Y = 8'b00111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 849,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110100; Y = 8'b01100110; // Expected: {'Z': -7752}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110100; Y = 8'b01100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 850,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7752
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110011; Y = 8'b10010011; // Expected: {'Z': 1417}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110011; Y = 8'b10010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 851,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1417
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110111; Y = 8'b10011111; // Expected: {'Z': 873}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110111; Y = 8'b10011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 852,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 873
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001100; Y = 8'b00111011; // Expected: {'Z': 708}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001100; Y = 8'b00111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 853,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 708
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000101; Y = 8'b11111010; // Expected: {'Z': -30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000101; Y = 8'b11111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 854,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000000; Y = 8'b10011010; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000000; Y = 8'b10011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 855,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000110; Y = 8'b01000111; // Expected: {'Z': -8662}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000110; Y = 8'b01000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 856,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8662
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011100; Y = 8'b00011011; // Expected: {'Z': -2700}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011100; Y = 8'b00011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 857,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000101; Y = 8'b00011000; // Expected: {'Z': 1656}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000101; Y = 8'b00011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 858,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1656
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110110; Y = 8'b01011011; // Expected: {'Z': 10738}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110110; Y = 8'b01011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 859,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10738
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010111; Y = 8'b10110000; // Expected: {'Z': 3280}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010111; Y = 8'b10110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 860,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010000; Y = 8'b01110110; // Expected: {'Z': 1888}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010000; Y = 8'b01110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 861,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001000; Y = 8'b00110101; // Expected: {'Z': 424}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001000; Y = 8'b00110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 862,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 424
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011100; Y = 8'b10000000; // Expected: {'Z': 4608}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011100; Y = 8'b10000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 863,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4608
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010111; Y = 8'b01011000; // Expected: {'Z': 2024}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010111; Y = 8'b01011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 864,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100010; Y = 8'b00110011; // Expected: {'Z': -4794}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100010; Y = 8'b00110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 865,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4794
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111001; Y = 8'b01011001; // Expected: {'Z': 5073}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111001; Y = 8'b01011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 866,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5073
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010000; Y = 8'b11011110; // Expected: {'Z': 1632}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010000; Y = 8'b11011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 867,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1632
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b10010111; // Expected: {'Z': -7140}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b10010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 868,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010010; Y = 8'b00010111; // Expected: {'Z': 1886}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010010; Y = 8'b00010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 869,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1886
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101000; Y = 8'b00101111; // Expected: {'Z': 1880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101000; Y = 8'b00101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 870,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111101; Y = 8'b01000100; // Expected: {'Z': -204}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111101; Y = 8'b01000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 871,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111000; Y = 8'b10101001; // Expected: {'Z': -10440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111000; Y = 8'b10101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 872,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101101; Y = 8'b01101010; // Expected: {'Z': 4770}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101101; Y = 8'b01101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 873,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4770
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100101; Y = 8'b10111000; // Expected: {'Z': 1944}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100101; Y = 8'b10111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 874,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011000; Y = 8'b01111011; // Expected: {'Z': 2952}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011000; Y = 8'b01111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 875,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2952
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000110; Y = 8'b11111000; // Expected: {'Z': -560}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000110; Y = 8'b11111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 876,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111111; Y = 8'b00000010; // Expected: {'Z': 254}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111111; Y = 8'b00000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 877,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110101; Y = 8'b01111101; // Expected: {'Z': -9375}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110101; Y = 8'b01111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 878,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9375
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101001; Y = 8'b00100101; // Expected: {'Z': -851}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101001; Y = 8'b00100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 879,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -851
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100110; Y = 8'b11000110; // Expected: {'Z': 1508}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100110; Y = 8'b11000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 880,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1508
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000110; Y = 8'b01011001; // Expected: {'Z': -5162}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000110; Y = 8'b01011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 881,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100111; Y = 8'b10010010; // Expected: {'Z': 9790}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100111; Y = 8'b10010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 882,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9790
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101111; Y = 8'b01111110; // Expected: {'Z': 13986}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101111; Y = 8'b01111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 883,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 13986
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001010; Y = 8'b01000010; // Expected: {'Z': -3564}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001010; Y = 8'b01000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 884,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3564
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110100; Y = 8'b10100101; // Expected: {'Z': 1092}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110100; Y = 8'b10100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 885,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1092
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110100; Y = 8'b10010101; // Expected: {'Z': 8132}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110100; Y = 8'b10010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 886,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110011; Y = 8'b00111100; // Expected: {'Z': -4620}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110011; Y = 8'b00111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 887,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000010; Y = 8'b01101011; // Expected: {'Z': -6634}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000010; Y = 8'b01101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 888,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6634
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001101; Y = 8'b01011110; // Expected: {'Z': -10810}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001101; Y = 8'b01011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 889,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10810
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010001; Y = 8'b00111110; // Expected: {'Z': 1054}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010001; Y = 8'b00111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 890,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1054
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100100; Y = 8'b01010000; // Expected: {'Z': 8000}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100100; Y = 8'b01010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 891,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010100; Y = 8'b00011101; // Expected: {'Z': 2436}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010100; Y = 8'b00011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 892,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2436
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101101; Y = 8'b00111001; // Expected: {'Z': -1083}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101101; Y = 8'b00111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 893,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1083
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100000; Y = 8'b00001000; // Expected: {'Z': 256}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100000; Y = 8'b00001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 894,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 256
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010111; Y = 8'b01011110; // Expected: {'Z': -3854}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010111; Y = 8'b01011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 895,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3854
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000011; Y = 8'b00010100; // Expected: {'Z': 1340}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000011; Y = 8'b00010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 896,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111000; Y = 8'b01011111; // Expected: {'Z': -760}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111000; Y = 8'b01011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 897,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110011; Y = 8'b10100101; // Expected: {'Z': -10465}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110011; Y = 8'b10100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 898,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10465
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111011; Y = 8'b10010100; // Expected: {'Z': 540}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111011; Y = 8'b10010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 899,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110011; Y = 8'b00111110; // Expected: {'Z': -4774}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110011; Y = 8'b00111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 900,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4774
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111001; Y = 8'b10110011; // Expected: {'Z': -4389}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111001; Y = 8'b10110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 901,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4389
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011110; Y = 8'b11101010; // Expected: {'Z': -2068}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011110; Y = 8'b11101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 902,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2068
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b00110011; // Expected: {'Z': 3774}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b00110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 903,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3774
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000001; Y = 8'b11110110; // Expected: {'Z': 630}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000001; Y = 8'b11110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 904,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 630
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b01111010; // Expected: {'Z': 8784}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b01111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 905,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111100; Y = 8'b11110000; // Expected: {'Z': 64}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111100; Y = 8'b11110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 906,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011110; Y = 8'b01000001; // Expected: {'Z': 1950}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011110; Y = 8'b01000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 907,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010110; Y = 8'b11001000; // Expected: {'Z': 5936}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010110; Y = 8'b11001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 908,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5936
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000000; Y = 8'b01010010; // Expected: {'Z': 5248}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000000; Y = 8'b01010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 909,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001101; Y = 8'b00111001; // Expected: {'Z': -6555}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001101; Y = 8'b00111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 910,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6555
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101010; Y = 8'b01011001; // Expected: {'Z': -1958}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101010; Y = 8'b01011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 911,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1958
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101110; Y = 8'b00001111; // Expected: {'Z': -270}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101110; Y = 8'b00001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 912,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -270
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010011; Y = 8'b00011010; // Expected: {'Z': -2834}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010011; Y = 8'b00011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 913,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2834
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010010; Y = 8'b11011001; // Expected: {'Z': -3198}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010010; Y = 8'b11011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 914,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b11111100; // Expected: {'Z': 328}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b11111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 915,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 328
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011101; Y = 8'b00101011; // Expected: {'Z': -4257}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011101; Y = 8'b00101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 916,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4257
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011111; Y = 8'b01100001; // Expected: {'Z': -3201}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011111; Y = 8'b01100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 917,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b10110110; // Expected: {'Z': -444}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b10110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 918,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -444
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010011; Y = 8'b01101100; // Expected: {'Z': -4860}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010011; Y = 8'b01101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 919,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4860
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101101; Y = 8'b10101000; // Expected: {'Z': -9592}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101101; Y = 8'b10101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 920,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9592
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010001; Y = 8'b01111000; // Expected: {'Z': 2040}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010001; Y = 8'b01111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 921,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011100; Y = 8'b01101001; // Expected: {'Z': 2940}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011100; Y = 8'b01101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 922,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2940
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101010; Y = 8'b10101100; // Expected: {'Z': -3528}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101010; Y = 8'b10101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 923,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111001; Y = 8'b01001000; // Expected: {'Z': 8712}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111001; Y = 8'b01001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 924,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8712
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001011; Y = 8'b01010101; // Expected: {'Z': -4505}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001011; Y = 8'b01010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 925,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4505
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110010; Y = 8'b10100110; // Expected: {'Z': 1260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110010; Y = 8'b10100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 926,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110110; Y = 8'b01011111; // Expected: {'Z': 11210}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110110; Y = 8'b01011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 927,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001100; Y = 8'b10100011; // Expected: {'Z': -7068}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001100; Y = 8'b10100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 928,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7068
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101110; Y = 8'b10010101; // Expected: {'Z': 1926}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101110; Y = 8'b10010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 929,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1926
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010100; Y = 8'b00101001; // Expected: {'Z': -1804}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010100; Y = 8'b00101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 930,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1804
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100110; Y = 8'b01011100; // Expected: {'Z': -8280}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100110; Y = 8'b01011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 931,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011010; Y = 8'b00110010; // Expected: {'Z': 1300}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011010; Y = 8'b00110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 932,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b01011101; // Expected: {'Z': 186}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b01011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 933,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b01111001; // Expected: {'Z': 8712}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b01111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 934,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8712
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000011; Y = 8'b11010011; // Expected: {'Z': -3015}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000011; Y = 8'b11010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 935,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3015
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100001; Y = 8'b10111011; // Expected: {'Z': -2277}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100001; Y = 8'b10111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 936,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2277
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b01001001; // Expected: {'Z': -6351}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b01001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 937,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6351
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111110; Y = 8'b00111110; // Expected: {'Z': 3844}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111110; Y = 8'b00111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 938,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3844
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101110; Y = 8'b11100101; // Expected: {'Z': 486}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101110; Y = 8'b11100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 939,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 486
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b01110111; // Expected: {'Z': 8092}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b01110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 940,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8092
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b10011100; // Expected: {'Z': -7200}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b10011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 941,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001100; Y = 8'b10100000; // Expected: {'Z': 4992}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001100; Y = 8'b10100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 942,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4992
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110001; Y = 8'b11111101; // Expected: {'Z': 237}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110001; Y = 8'b11111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 943,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 237
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000111; Y = 8'b10100011; // Expected: {'Z': -6603}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000111; Y = 8'b10100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 944,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6603
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010000; Y = 8'b01110010; // Expected: {'Z': 1824}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010000; Y = 8'b01110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 945,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1824
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110011; Y = 8'b11101100; // Expected: {'Z': -1020}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110011; Y = 8'b11101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 946,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1020
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010010; Y = 8'b01101101; // Expected: {'Z': 8938}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010010; Y = 8'b01101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 947,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8938
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010011; Y = 8'b11101100; // Expected: {'Z': 900}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010011; Y = 8'b11101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 948,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101011; Y = 8'b00111101; // Expected: {'Z': 6527}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101011; Y = 8'b00111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 949,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6527
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100101; Y = 8'b11001010; // Expected: {'Z': -5454}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100101; Y = 8'b11001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 950,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5454
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101101; Y = 8'b01000011; // Expected: {'Z': -5561}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101101; Y = 8'b01000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 951,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5561
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b01011011; // Expected: {'Z': 6734}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b01011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 952,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6734
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000011; Y = 8'b00111011; // Expected: {'Z': 3953}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000011; Y = 8'b00111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 953,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3953
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b11000010; // Expected: {'Z': 5394}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b11000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 954,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5394
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010010; Y = 8'b00000100; // Expected: {'Z': -440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010010; Y = 8'b00000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 955,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101111; Y = 8'b00110110; // Expected: {'Z': 5994}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101111; Y = 8'b00110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 956,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5994
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100001; Y = 8'b10110001; // Expected: {'Z': 7505}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100001; Y = 8'b10110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 957,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7505
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101101; Y = 8'b01001010; // Expected: {'Z': -1406}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101101; Y = 8'b01001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 958,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1406
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000101; Y = 8'b01111100; // Expected: {'Z': 8556}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000101; Y = 8'b01111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 959,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8556
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100101; Y = 8'b11001101; // Expected: {'Z': 1377}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100101; Y = 8'b11001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 960,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1377
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000101; Y = 8'b01001000; // Expected: {'Z': 360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000101; Y = 8'b01001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 961,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101110; Y = 8'b10001101; // Expected: {'Z': 2070}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101110; Y = 8'b10001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 962,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2070
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000111; Y = 8'b01011110; // Expected: {'Z': 658}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000111; Y = 8'b01011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 963,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 658
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b01101010; // Expected: {'Z': 4982}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b01101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 964,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4982
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011001; Y = 8'b10001110; // Expected: {'Z': 4446}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011001; Y = 8'b10001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 965,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4446
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101010; Y = 8'b11110100; // Expected: {'Z': 1032}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101010; Y = 8'b11110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 966,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1032
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100100; Y = 8'b00010100; // Expected: {'Z': 2000}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100100; Y = 8'b00010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 967,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101011; Y = 8'b00101111; // Expected: {'Z': 5029}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101011; Y = 8'b00101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 968,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5029
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b01110110; // Expected: {'Z': -9912}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b01110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 969,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9912
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011100; Y = 8'b00000011; // Expected: {'Z': -300}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011100; Y = 8'b00000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 970,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b00011000; // Expected: {'Z': 2472}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b00011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 971,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2472
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011110; Y = 8'b00010110; // Expected: {'Z': 660}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011110; Y = 8'b00010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 972,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111111; Y = 8'b10011001; // Expected: {'Z': 6695}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111111; Y = 8'b10011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 973,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6695
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111101; Y = 8'b10100011; // Expected: {'Z': -11625}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111101; Y = 8'b10100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 974,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11625
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010100; Y = 8'b00100100; // Expected: {'Z': -1584}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010100; Y = 8'b00100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 975,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1584
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010111; Y = 8'b10010101; // Expected: {'Z': 4387}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010111; Y = 8'b10010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 976,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4387
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011010; Y = 8'b11100000; // Expected: {'Z': -2880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011010; Y = 8'b11100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 977,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111111; Y = 8'b11010110; // Expected: {'Z': -5334}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111111; Y = 8'b11010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 978,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5334
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100110; Y = 8'b10001011; // Expected: {'Z': 3042}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100110; Y = 8'b10001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 979,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3042
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011110; Y = 8'b11000011; // Expected: {'Z': -1830}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011110; Y = 8'b11000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 980,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1830
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111010; Y = 8'b11100110; // Expected: {'Z': -3172}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111010; Y = 8'b11100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 981,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110010; Y = 8'b01110110; // Expected: {'Z': -1652}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110010; Y = 8'b01110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 982,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1652
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001110; Y = 8'b11010111; // Expected: {'Z': -574}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001110; Y = 8'b11010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 983,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -574
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100110; Y = 8'b10100100; // Expected: {'Z': 8280}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100110; Y = 8'b10100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 984,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111011; Y = 8'b00100111; // Expected: {'Z': -195}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111011; Y = 8'b00100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 985,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101100; Y = 8'b00111000; // Expected: {'Z': -1120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101100; Y = 8'b00111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 986,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110100; Y = 8'b01010110; // Expected: {'Z': 4472}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110100; Y = 8'b01010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 987,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4472
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010010; Y = 8'b01111001; // Expected: {'Z': 2178}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010010; Y = 8'b01111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 988,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111001; Y = 8'b10000100; // Expected: {'Z': 8804}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111001; Y = 8'b10000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 989,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8804
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011100; Y = 8'b10001110; // Expected: {'Z': -3192}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011100; Y = 8'b10001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 990,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111111; Y = 8'b11001000; // Expected: {'Z': 3640}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111111; Y = 8'b11001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 991,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100001; Y = 8'b01011100; // Expected: {'Z': 8924}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100001; Y = 8'b01011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 992,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8924
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000010; Y = 8'b10011011; // Expected: {'Z': 6262}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000010; Y = 8'b10011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 993,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6262
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001001; Y = 8'b01101100; // Expected: {'Z': -5940}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001001; Y = 8'b01101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 994,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5940
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011000; Y = 8'b01100101; // Expected: {'Z': -4040}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011000; Y = 8'b01100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 995,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b01001000; // Expected: {'Z': 1080}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b01001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 996,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b01101011; // Expected: {'Z': -11877}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b01101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 997,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11877
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011111; Y = 8'b00101011; // Expected: {'Z': -4171}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011111; Y = 8'b00101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 998,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110101; Y = 8'b10011010; // Expected: {'Z': 1122}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110101; Y = 8'b10011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 999,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b00100000; // Expected: {'Z': -896}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b00100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1000,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b10111010; // Expected: {'Z': -8610}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b10111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1001,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8610
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011010; Y = 8'b10110101; // Expected: {'Z': -6750}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011010; Y = 8'b10110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1002,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100010; Y = 8'b11011101; // Expected: {'Z': 3290}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100010; Y = 8'b11011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1003,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3290
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010111; Y = 8'b01111011; // Expected: {'Z': 2829}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010111; Y = 8'b01111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1004,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2829
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101010; Y = 8'b10100101; // Expected: {'Z': 2002}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101010; Y = 8'b10100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1005,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2002
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110111; Y = 8'b10000100; // Expected: {'Z': 9052}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110111; Y = 8'b10000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1006,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9052
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b10011000; // Expected: {'Z': -4056}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b10011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1007,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4056
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001001; Y = 8'b01101001; // Expected: {'Z': 7665}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001001; Y = 8'b01101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1008,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7665
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111001; Y = 8'b11001101; // Expected: {'Z': 357}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111001; Y = 8'b11001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1009,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 357
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000110; Y = 8'b10111100; // Expected: {'Z': 3944}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000110; Y = 8'b10111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1010,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001100; Y = 8'b10101011; // Expected: {'Z': -6460}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001100; Y = 8'b10101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1011,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6460
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111001; Y = 8'b00000011; // Expected: {'Z': -213}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111001; Y = 8'b00000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1012,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b00111100; // Expected: {'Z': -6660}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b00111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1013,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001011; Y = 8'b01111010; // Expected: {'Z': -14274}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001011; Y = 8'b01111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1014,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -14274
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000111; Y = 8'b01101010; // Expected: {'Z': -6042}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000111; Y = 8'b01101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1015,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6042
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110010; Y = 8'b01010010; // Expected: {'Z': -6396}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110010; Y = 8'b01010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1016,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6396
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010100; Y = 8'b00101001; // Expected: {'Z': -4428}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010100; Y = 8'b00101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1017,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4428
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b01011011; // Expected: {'Z': -2548}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b01011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1018,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2548
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b11010111; // Expected: {'Z': -4592}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b11010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1019,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4592
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b11011010; // Expected: {'Z': -76}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b11011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1020,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010110; Y = 8'b01010110; // Expected: {'Z': 7396}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010110; Y = 8'b01010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1021,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7396
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100010; Y = 8'b01010110; // Expected: {'Z': -2580}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100010; Y = 8'b01010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1022,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111011; Y = 8'b01110100; // Expected: {'Z': -580}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111011; Y = 8'b01110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1023,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001011; Y = 8'b01100001; // Expected: {'Z': 7275}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001011; Y = 8'b01100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1024,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7275
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b11011001; // Expected: {'Z': -2379}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b11011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1025,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2379
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000000; Y = 8'b11010010; // Expected: {'Z': 2944}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000000; Y = 8'b11010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1026,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b10110001; // Expected: {'Z': 6873}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b10110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1027,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6873
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111111; Y = 8'b10100101; // Expected: {'Z': -5733}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111111; Y = 8'b10100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1028,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5733
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001011; Y = 8'b11111001; // Expected: {'Z': 819}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001011; Y = 8'b11111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1029,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 819
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100110; Y = 8'b10000001; // Expected: {'Z': 11430}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100110; Y = 8'b10000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1030,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000011; Y = 8'b01000010; // Expected: {'Z': -4026}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000011; Y = 8'b01000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1031,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4026
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000010; Y = 8'b01111111; // Expected: {'Z': 8382}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000010; Y = 8'b01111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1032,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8382
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b11111111; // Expected: {'Z': -96}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b11111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1033,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011110; Y = 8'b00001111; // Expected: {'Z': -1470}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011110; Y = 8'b00001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1034,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1470
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011110; Y = 8'b00100110; // Expected: {'Z': 3572}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011110; Y = 8'b00100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1035,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3572
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100010; Y = 8'b10100100; // Expected: {'Z': 8648}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100010; Y = 8'b10100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1036,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010010; Y = 8'b11010001; // Expected: {'Z': 2162}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010010; Y = 8'b11010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1037,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100110; Y = 8'b00101000; // Expected: {'Z': 4080}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100110; Y = 8'b00101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1038,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101001; Y = 8'b10110101; // Expected: {'Z': -7875}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101001; Y = 8'b10110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1039,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7875
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b11001111; // Expected: {'Z': -4312}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b11001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1040,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4312
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110011; Y = 8'b00011101; // Expected: {'Z': 3335}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110011; Y = 8'b00011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1041,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3335
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100000; Y = 8'b00000101; // Expected: {'Z': -160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100000; Y = 8'b00000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1042,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011111; Y = 8'b00101001; // Expected: {'Z': -3977}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011111; Y = 8'b00101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1043,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3977
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b10011100; // Expected: {'Z': -200}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b10011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1044,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001001; Y = 8'b10100110; // Expected: {'Z': 4950}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001001; Y = 8'b10100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1045,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110011; Y = 8'b11010011; // Expected: {'Z': 3465}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110011; Y = 8'b11010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1046,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3465
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111001; Y = 8'b01111001; // Expected: {'Z': 14641}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111001; Y = 8'b01111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1047,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 14641
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110111; Y = 8'b10110010; // Expected: {'Z': 702}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110111; Y = 8'b10110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1048,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 702
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001101; Y = 8'b10100000; // Expected: {'Z': -7392}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001101; Y = 8'b10100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1049,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100011; Y = 8'b10010110; // Expected: {'Z': 3074}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100011; Y = 8'b10010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1050,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3074
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010111; Y = 8'b11011111; // Expected: {'Z': -2871}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010111; Y = 8'b11011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1051,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2871
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111010; Y = 8'b10101100; // Expected: {'Z': 504}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111010; Y = 8'b10101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1052,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111101; Y = 8'b10001100; // Expected: {'Z': 7772}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111101; Y = 8'b10001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1053,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7772
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000011; Y = 8'b11100100; // Expected: {'Z': 1708}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000011; Y = 8'b11100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1054,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1708
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111010; Y = 8'b10011110; // Expected: {'Z': -5684}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111010; Y = 8'b10011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1055,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5684
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100001; Y = 8'b00001010; // Expected: {'Z': 970}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100001; Y = 8'b00001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1056,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 970
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b00101111; // Expected: {'Z': 2538}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b00101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1057,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2538
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b11100011; // Expected: {'Z': 1624}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b11100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1058,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b00001100; // Expected: {'Z': 348}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b00001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1059,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 348
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110001; Y = 8'b01011110; // Expected: {'Z': -1410}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110001; Y = 8'b01011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1060,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1410
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101000; Y = 8'b10100100; // Expected: {'Z': 8096}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101000; Y = 8'b10100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1061,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8096
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100001; Y = 8'b10001101; // Expected: {'Z': -3795}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100001; Y = 8'b10001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1062,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3795
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010111; Y = 8'b01101011; // Expected: {'Z': 2461}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010111; Y = 8'b01101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1063,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2461
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100100; Y = 8'b01000000; // Expected: {'Z': -5888}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100100; Y = 8'b01000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1064,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111010; Y = 8'b11000110; // Expected: {'Z': 4060}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111010; Y = 8'b11000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1065,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101011; Y = 8'b10101101; // Expected: {'Z': 1743}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101011; Y = 8'b10101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1066,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1743
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000001; Y = 8'b00111110; // Expected: {'Z': -7874}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000001; Y = 8'b00111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1067,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7874
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100111; Y = 8'b11100001; // Expected: {'Z': 2759}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100111; Y = 8'b11100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1068,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2759
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100011; Y = 8'b11010011; // Expected: {'Z': 4185}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100011; Y = 8'b11010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1069,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111010; Y = 8'b10001000; // Expected: {'Z': 8400}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111010; Y = 8'b10001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1070,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011001; Y = 8'b00111110; // Expected: {'Z': 5518}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011001; Y = 8'b00111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1071,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5518
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b01011101; // Expected: {'Z': -4743}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b01011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1072,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4743
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100111; Y = 8'b01000010; // Expected: {'Z': -1650}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100111; Y = 8'b01000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1073,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b00011000; // Expected: {'Z': 1728}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b00011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1074,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110111; Y = 8'b10111011; // Expected: {'Z': 621}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110111; Y = 8'b10111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1075,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 621
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b10110111; // Expected: {'Z': -1387}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b10110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1076,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1387
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111111; Y = 8'b00100100; // Expected: {'Z': 2268}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111111; Y = 8'b00100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1077,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2268
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111011; Y = 8'b01110100; // Expected: {'Z': 6844}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111011; Y = 8'b01110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1078,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6844
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011101; Y = 8'b11011110; // Expected: {'Z': 1190}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011101; Y = 8'b11011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1079,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110100; Y = 8'b11101010; // Expected: {'Z': 1672}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110100; Y = 8'b11101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1080,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111010; Y = 8'b00111001; // Expected: {'Z': -342}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111010; Y = 8'b00111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1081,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -342
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001011; Y = 8'b11011101; // Expected: {'Z': -385}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001011; Y = 8'b11011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1082,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -385
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110100; Y = 8'b00101011; // Expected: {'Z': -516}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110100; Y = 8'b00101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1083,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -516
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001101; Y = 8'b00010010; // Expected: {'Z': 1386}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001101; Y = 8'b00010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1084,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1386
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110010; Y = 8'b11001011; // Expected: {'Z': -2650}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110010; Y = 8'b11001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1085,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010111; Y = 8'b01100101; // Expected: {'Z': -10605}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010111; Y = 8'b01100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1086,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10605
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001111; Y = 8'b10110001; // Expected: {'Z': 3871}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001111; Y = 8'b10110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1087,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3871
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101000; Y = 8'b11110101; // Expected: {'Z': -440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101000; Y = 8'b11110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1088,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011110; Y = 8'b11011001; // Expected: {'Z': -3666}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011110; Y = 8'b11011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1089,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3666
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010001; Y = 8'b01100010; // Expected: {'Z': 1666}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010001; Y = 8'b01100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1090,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1666
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101000; Y = 8'b01011110; // Expected: {'Z': -2256}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101000; Y = 8'b01011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1091,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2256
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111001; Y = 8'b01010110; // Expected: {'Z': -6106}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111001; Y = 8'b01010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1092,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000100; Y = 8'b01000111; // Expected: {'Z': -4260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000100; Y = 8'b01000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1093,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010111; Y = 8'b10001000; // Expected: {'Z': -2760}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010111; Y = 8'b10001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1094,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111110; Y = 8'b00101111; // Expected: {'Z': 2914}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111110; Y = 8'b00101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1095,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2914
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111111; Y = 8'b11011111; // Expected: {'Z': -2079}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111111; Y = 8'b11011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1096,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2079
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011111; Y = 8'b01111011; // Expected: {'Z': 11685}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011111; Y = 8'b01111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1097,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11685
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010010; Y = 8'b01001010; // Expected: {'Z': -3404}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010010; Y = 8'b01001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1098,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3404
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001011; Y = 8'b00001000; // Expected: {'Z': 600}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001011; Y = 8'b00001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1099,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b01100000; // Expected: {'Z': 4512}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b01100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1100,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4512
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110011; Y = 8'b10111100; // Expected: {'Z': -7820}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110011; Y = 8'b10111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1101,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b00111000; // Expected: {'Z': 1064}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b00111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1102,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1064
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011011; Y = 8'b10000101; // Expected: {'Z': 12423}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011011; Y = 8'b10000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1103,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 12423
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010011; Y = 8'b01101000; // Expected: {'Z': 8632}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010011; Y = 8'b01101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1104,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8632
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000111; Y = 8'b00011111; // Expected: {'Z': -1767}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000111; Y = 8'b00011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1105,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1767
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010111; Y = 8'b00101001; // Expected: {'Z': -1681}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010111; Y = 8'b00101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1106,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1681
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010000; Y = 8'b00011101; // Expected: {'Z': -1392}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010000; Y = 8'b00011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1107,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101001; Y = 8'b10000100; // Expected: {'Z': -13020}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101001; Y = 8'b10000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1108,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -13020
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011010; Y = 8'b10010111; // Expected: {'Z': -9450}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011010; Y = 8'b10010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1109,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010111; Y = 8'b10111111; // Expected: {'Z': -5655}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010111; Y = 8'b10111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1110,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5655
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111100; Y = 8'b11111001; // Expected: {'Z': -868}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111100; Y = 8'b11111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1111,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -868
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110111; Y = 8'b00100111; // Expected: {'Z': 4641}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110111; Y = 8'b00100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1112,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4641
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b01001110; // Expected: {'Z': 5304}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b01001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1113,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5304
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001111; Y = 8'b11111001; // Expected: {'Z': 343}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001111; Y = 8'b11111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1114,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 343
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100010; Y = 8'b01100001; // Expected: {'Z': -2910}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100010; Y = 8'b01100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1115,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2910
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010001; Y = 8'b10100001; // Expected: {'Z': 4465}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010001; Y = 8'b10100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1116,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4465
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111101; Y = 8'b01001010; // Expected: {'Z': -4958}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111101; Y = 8'b01001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1117,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4958
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111110; Y = 8'b01111000; // Expected: {'Z': -240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111110; Y = 8'b01111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1118,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010000; Y = 8'b01001001; // Expected: {'Z': -3504}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010000; Y = 8'b01001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1119,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011111; Y = 8'b00101010; // Expected: {'Z': 3990}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011111; Y = 8'b00101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1120,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3990
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101101; Y = 8'b10000100; // Expected: {'Z': -13516}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101101; Y = 8'b10000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1121,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -13516
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111010; Y = 8'b11101101; // Expected: {'Z': 1330}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111010; Y = 8'b11101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1122,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1330
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100000; Y = 8'b00001011; // Expected: {'Z': 352}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100000; Y = 8'b00001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1123,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110001; Y = 8'b10111000; // Expected: {'Z': 5688}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110001; Y = 8'b10111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1124,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5688
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100010; Y = 8'b00100111; // Expected: {'Z': 1326}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100010; Y = 8'b00100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1125,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1326
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110110; Y = 8'b00011100; // Expected: {'Z': -2072}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110110; Y = 8'b00011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1126,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2072
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000000; Y = 8'b10101100; // Expected: {'Z': -5376}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000000; Y = 8'b10101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1127,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5376
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b00000001; // Expected: {'Z': -68}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b00000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1128,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111011; Y = 8'b11111011; // Expected: {'Z': 345}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111011; Y = 8'b11111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1129,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 345
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111011; Y = 8'b01010010; // Expected: {'Z': 4838}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111011; Y = 8'b01010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1130,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4838
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001111; Y = 8'b00110001; // Expected: {'Z': 3871}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001111; Y = 8'b00110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1131,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3871
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001000; Y = 8'b10111110; // Expected: {'Z': -528}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001000; Y = 8'b10111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1132,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b11000111; // Expected: {'Z': -855}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b11000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1133,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -855
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000001; Y = 8'b00110001; // Expected: {'Z': 3185}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000001; Y = 8'b00110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1134,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b00000110; // Expected: {'Z': 54}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b00000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1135,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000110; Y = 8'b00100010; // Expected: {'Z': -4148}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000110; Y = 8'b00100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1136,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111111; Y = 8'b00000001; // Expected: {'Z': -1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111111; Y = 8'b00000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1137,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001110; Y = 8'b11001011; // Expected: {'Z': -4134}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001110; Y = 8'b11001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1138,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000101; Y = 8'b11011011; // Expected: {'Z': 4551}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000101; Y = 8'b11011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1139,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4551
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101110; Y = 8'b11000101; // Expected: {'Z': -6490}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101110; Y = 8'b11000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1140,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6490
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011010; Y = 8'b01101110; // Expected: {'Z': -11220}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011010; Y = 8'b01101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1141,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100111; Y = 8'b11010001; // Expected: {'Z': 1175}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100111; Y = 8'b11010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1142,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100101; Y = 8'b01001010; // Expected: {'Z': 7474}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100101; Y = 8'b01001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1143,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7474
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100001; Y = 8'b00111100; // Expected: {'Z': -1860}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100001; Y = 8'b00111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1144,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1860
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110100; Y = 8'b01001100; // Expected: {'Z': 8816}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110100; Y = 8'b01001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1145,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011011; Y = 8'b11010101; // Expected: {'Z': 4343}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011011; Y = 8'b11010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1146,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4343
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011110; Y = 8'b01111000; // Expected: {'Z': 11280}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011110; Y = 8'b01111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1147,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111000; Y = 8'b00110110; // Expected: {'Z': 3024}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111000; Y = 8'b00110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1148,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b11100101; // Expected: {'Z': -2592}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b11100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1149,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2592
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011001; Y = 8'b00111100; // Expected: {'Z': -6180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011001; Y = 8'b00111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1150,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110001; Y = 8'b01111111; // Expected: {'Z': -10033}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110001; Y = 8'b01111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1151,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10033
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001111; Y = 8'b11001010; // Expected: {'Z': 2646}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001111; Y = 8'b11001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1152,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2646
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111111; Y = 8'b00101101; // Expected: {'Z': 2835}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111111; Y = 8'b00101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1153,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2835
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010010; Y = 8'b10110011; // Expected: {'Z': -1386}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010010; Y = 8'b10110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1154,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1386
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000011; Y = 8'b10001010; // Expected: {'Z': 14750}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000011; Y = 8'b10001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1155,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 14750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000110; Y = 8'b11101100; // Expected: {'Z': 1160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000110; Y = 8'b11101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1156,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011110; Y = 8'b11100010; // Expected: {'Z': -2820}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011110; Y = 8'b11100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1157,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101001; Y = 8'b01000001; // Expected: {'Z': -1495}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101001; Y = 8'b01000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1158,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1495
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110010; Y = 8'b10110101; // Expected: {'Z': -8550}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110010; Y = 8'b10110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1159,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010001; Y = 8'b10111100; // Expected: {'Z': -1156}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010001; Y = 8'b10111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1160,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000001; Y = 8'b00111101; // Expected: {'Z': 61}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000001; Y = 8'b00111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1161,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011011; Y = 8'b00100011; // Expected: {'Z': 3185}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011011; Y = 8'b00100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1162,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b01010010; // Expected: {'Z': 9184}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b01010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1163,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b11000100; // Expected: {'Z': -2640}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b11000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1164,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000010; Y = 8'b01101011; // Expected: {'Z': 7062}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000010; Y = 8'b01101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1165,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7062
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100110; Y = 8'b01000011; // Expected: {'Z': 2546}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100110; Y = 8'b01000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1166,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001101; Y = 8'b00110101; // Expected: {'Z': -6095}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001101; Y = 8'b00110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1167,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6095
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101000; Y = 8'b01110111; // Expected: {'Z': 4760}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101000; Y = 8'b01110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1168,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110010; Y = 8'b10110010; // Expected: {'Z': -3900}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110010; Y = 8'b10110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1169,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000000; Y = 8'b10011011; // Expected: {'Z': 12928}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000000; Y = 8'b10011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1170,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 12928
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100010; Y = 8'b01011100; // Expected: {'Z': -2760}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100010; Y = 8'b01011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1171,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b11000001; // Expected: {'Z': 5481}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b11000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1172,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5481
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001110; Y = 8'b10001100; // Expected: {'Z': 13224}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001110; Y = 8'b10001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1173,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 13224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001110; Y = 8'b10111010; // Expected: {'Z': 3500}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001110; Y = 8'b10111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1174,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100001; Y = 8'b00101000; // Expected: {'Z': -3800}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100001; Y = 8'b00101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1175,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011110; Y = 8'b11010110; // Expected: {'Z': -1260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011110; Y = 8'b11010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1176,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011000; Y = 8'b01101110; // Expected: {'Z': 2640}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011000; Y = 8'b01101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1177,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011011; Y = 8'b11001110; // Expected: {'Z': 5050}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011011; Y = 8'b11001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1178,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110011; Y = 8'b11000100; // Expected: {'Z': -3060}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110011; Y = 8'b11000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1179,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001010; Y = 8'b01000100; // Expected: {'Z': -3672}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001010; Y = 8'b01000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1180,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b11000110; // Expected: {'Z': -116}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b11000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1181,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110110; Y = 8'b10110011; // Expected: {'Z': 770}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110110; Y = 8'b10110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1182,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 770
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101100; Y = 8'b00101010; // Expected: {'Z': 4536}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101100; Y = 8'b00101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1183,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4536
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b01011000; // Expected: {'Z': -2464}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b01011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1184,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001010; Y = 8'b00010100; // Expected: {'Z': -2360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001010; Y = 8'b00010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1185,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010000; Y = 8'b11101101; // Expected: {'Z': 2128}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010000; Y = 8'b11101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1186,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000000; Y = 8'b11101001; // Expected: {'Z': 2944}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000000; Y = 8'b11101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1187,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110110; Y = 8'b11100000; // Expected: {'Z': 320}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110110; Y = 8'b11100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1188,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111001; Y = 8'b00101011; // Expected: {'Z': -3053}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111001; Y = 8'b00101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1189,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3053
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010010; Y = 8'b00110101; // Expected: {'Z': -2438}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010010; Y = 8'b00110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1190,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2438
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110100; Y = 8'b10011111; // Expected: {'Z': 7372}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110100; Y = 8'b10011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1191,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7372
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b11011100; // Expected: {'Z': 1836}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b11011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1192,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1836
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b11010100; // Expected: {'Z': 3696}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b11010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1193,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3696
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000100; Y = 8'b11001101; // Expected: {'Z': 3060}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000100; Y = 8'b11001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1194,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001011; Y = 8'b01011011; // Expected: {'Z': 1001}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001011; Y = 8'b01011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1195,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1001
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000101; Y = 8'b11111011; // Expected: {'Z': -25}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000101; Y = 8'b11111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1196,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b00011000; // Expected: {'Z': 1632}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b00011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1197,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1632
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100110; Y = 8'b00101010; // Expected: {'Z': -1092}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100110; Y = 8'b00101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1198,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1092
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010001; Y = 8'b11111101; // Expected: {'Z': 141}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010001; Y = 8'b11111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1199,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111111; Y = 8'b11101110; // Expected: {'Z': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111111; Y = 8'b11101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1200,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010000; Y = 8'b01100000; // Expected: {'Z': -10752}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010000; Y = 8'b01100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1201,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10752
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100011; Y = 8'b01001000; // Expected: {'Z': -6696}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100011; Y = 8'b01001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1202,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6696
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000001; Y = 8'b11100010; // Expected: {'Z': -1950}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000001; Y = 8'b11100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1203,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000011; Y = 8'b10110000; // Expected: {'Z': 10000}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000011; Y = 8'b10110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1204,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100110; Y = 8'b00110101; // Expected: {'Z': -4770}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100110; Y = 8'b00110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1205,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4770
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111110; Y = 8'b11011110; // Expected: {'Z': -2108}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111110; Y = 8'b11011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1206,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011111; Y = 8'b00110011; // Expected: {'Z': -1683}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011111; Y = 8'b00110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1207,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1683
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110100; Y = 8'b00011011; // Expected: {'Z': -2052}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110100; Y = 8'b00011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1208,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2052
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001001; Y = 8'b00011001; // Expected: {'Z': -2975}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001001; Y = 8'b00011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1209,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2975
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000111; Y = 8'b11000101; // Expected: {'Z': -413}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000111; Y = 8'b11000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1210,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -413
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000100; Y = 8'b01111110; // Expected: {'Z': -15624}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000100; Y = 8'b01111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1211,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -15624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b10100111; // Expected: {'Z': -801}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b10100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1212,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -801
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b11000110; // Expected: {'Z': -5974}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b11000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1213,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5974
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010000; Y = 8'b01011100; // Expected: {'Z': 1472}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010000; Y = 8'b01011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1214,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1472
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b01010000; // Expected: {'Z': 1040}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b01010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1215,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101010; Y = 8'b10011001; // Expected: {'Z': 2266}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101010; Y = 8'b10011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1216,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2266
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b01000111; // Expected: {'Z': -5822}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b01000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1217,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5822
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b01011101; // Expected: {'Z': 5022}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b01011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1218,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5022
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000010; Y = 8'b11111110; // Expected: {'Z': 124}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000010; Y = 8'b11111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1219,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011101; Y = 8'b01011011; // Expected: {'Z': 8463}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011101; Y = 8'b01011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1220,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8463
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110000; Y = 8'b11001111; // Expected: {'Z': 784}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110000; Y = 8'b11001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1221,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001011; Y = 8'b11110010; // Expected: {'Z': -154}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001011; Y = 8'b11110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1222,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011001; Y = 8'b00110111; // Expected: {'Z': -5665}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011001; Y = 8'b00110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1223,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5665
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b11101001; // Expected: {'Z': 644}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b11101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1224,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 644
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111101; Y = 8'b11010000; // Expected: {'Z': -6000}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111101; Y = 8'b11010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1225,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010111; Y = 8'b00011100; // Expected: {'Z': 2436}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010111; Y = 8'b00011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1226,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2436
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b11111101; // Expected: {'Z': -63}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b11111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1227,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b01000100; // Expected: {'Z': -4624}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b01000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1228,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100001; Y = 8'b11011001; // Expected: {'Z': 3705}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100001; Y = 8'b11011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1229,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3705
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b11101101; // Expected: {'Z': 969}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b11101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1230,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 969
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001011; Y = 8'b11000001; // Expected: {'Z': -693}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001011; Y = 8'b11000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1231,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -693
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b10000011; // Expected: {'Z': -1875}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b10000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1232,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1875
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101101; Y = 8'b01000100; // Expected: {'Z': 3060}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101101; Y = 8'b01000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1233,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000001; Y = 8'b00000001; // Expected: {'Z': 65}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000001; Y = 8'b00000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1234,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001010; Y = 8'b10001001; // Expected: {'Z': 14042}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001010; Y = 8'b10001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1235,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 14042
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100010; Y = 8'b00000010; // Expected: {'Z': 68}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100010; Y = 8'b00000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1236,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111010; Y = 8'b00110000; // Expected: {'Z': -3360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111010; Y = 8'b00110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1237,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111100; Y = 8'b10011110; // Expected: {'Z': -12152}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111100; Y = 8'b10011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1238,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110000; Y = 8'b00001011; // Expected: {'Z': -880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110000; Y = 8'b00001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1239,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100000; Y = 8'b10101010; // Expected: {'Z': 2752}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100000; Y = 8'b10101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1240,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2752
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101101; Y = 8'b01000010; // Expected: {'Z': -1254}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101101; Y = 8'b01000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1241,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b10000011; // Expected: {'Z': -2625}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b10000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1242,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2625
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110111; Y = 8'b11001110; // Expected: {'Z': -5950}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110111; Y = 8'b11001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1243,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011010; Y = 8'b00101011; // Expected: {'Z': -4386}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011010; Y = 8'b00101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1244,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4386
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001001; Y = 8'b01110001; // Expected: {'Z': 8249}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001001; Y = 8'b01110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1245,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011001; Y = 8'b00111001; // Expected: {'Z': 5073}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011001; Y = 8'b00111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1246,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5073
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000011; Y = 8'b11101000; // Expected: {'Z': 3000}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000011; Y = 8'b11101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1247,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110010; Y = 8'b01011000; // Expected: {'Z': -1232}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110010; Y = 8'b01011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1248,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000100; Y = 8'b10100011; // Expected: {'Z': 5580}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000100; Y = 8'b10100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1249,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101000; Y = 8'b10011000; // Expected: {'Z': 9152}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101000; Y = 8'b10011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1250,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b10110101; // Expected: {'Z': -2700}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b10110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1251,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101011; Y = 8'b00100011; // Expected: {'Z': -735}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101011; Y = 8'b00100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1252,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -735
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011111; Y = 8'b00000010; // Expected: {'Z': 62}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011111; Y = 8'b00000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1253,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b01000000; // Expected: {'Z': -7104}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b01000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1254,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b00000110; // Expected: {'Z': -504}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b00000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1255,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011100; Y = 8'b10011010; // Expected: {'Z': 3672}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011100; Y = 8'b10011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1256,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100110; Y = 8'b01110001; // Expected: {'Z': 11526}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100110; Y = 8'b01110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1257,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11526
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110101; Y = 8'b00101111; // Expected: {'Z': 5499}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110101; Y = 8'b00101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1258,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5499
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010110; Y = 8'b00011110; // Expected: {'Z': -3180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010110; Y = 8'b00011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1259,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001110; Y = 8'b00101111; // Expected: {'Z': 3666}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001110; Y = 8'b00101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1260,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3666
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010010; Y = 8'b01110111; // Expected: {'Z': -5474}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010010; Y = 8'b01110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1261,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5474
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b11010011; // Expected: {'Z': -990}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b11010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1262,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -990
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100101; Y = 8'b00010011; // Expected: {'Z': -513}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100101; Y = 8'b00010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1263,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -513
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000011; Y = 8'b00001011; // Expected: {'Z': 737}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000011; Y = 8'b00001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1264,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 737
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100101; Y = 8'b00001110; // Expected: {'Z': 1414}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100101; Y = 8'b00001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1265,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1414
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010011; Y = 8'b11011010; // Expected: {'Z': -3154}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010011; Y = 8'b11011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1266,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100111; Y = 8'b10111101; // Expected: {'Z': 1675}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100111; Y = 8'b10111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1267,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1675
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101010; Y = 8'b01101111; // Expected: {'Z': -2442}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101010; Y = 8'b01101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1268,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2442
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b01001000; // Expected: {'Z': 432}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b01001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1269,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010001; Y = 8'b11101100; // Expected: {'Z': 940}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010001; Y = 8'b11101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1270,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 940
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100011; Y = 8'b00011101; // Expected: {'Z': -2697}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100011; Y = 8'b00011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1271,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2697
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100110; Y = 8'b11001000; // Expected: {'Z': -5712}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100110; Y = 8'b11001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1272,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5712
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b00101110; // Expected: {'Z': 414}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b00101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1273,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 414
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100110; Y = 8'b01111100; // Expected: {'Z': -3224}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100110; Y = 8'b01111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1274,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111000; Y = 8'b01000001; // Expected: {'Z': -520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111000; Y = 8'b01000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1275,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b00010100; // Expected: {'Z': 580}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b00010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1276,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100110; Y = 8'b11011010; // Expected: {'Z': 988}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100110; Y = 8'b11011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1277,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 988
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110100; Y = 8'b01010001; // Expected: {'Z': 9396}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110100; Y = 8'b01010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1278,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9396
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b01010101; // Expected: {'Z': 1615}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b01010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1279,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1615
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010110; Y = 8'b10101101; // Expected: {'Z': 3486}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010110; Y = 8'b10101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1280,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3486
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010100; Y = 8'b00111010; // Expected: {'Z': 1160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010100; Y = 8'b00111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1281,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111100; Y = 8'b10011010; // Expected: {'Z': 408}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111100; Y = 8'b10011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1282,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011011; Y = 8'b10100010; // Expected: {'Z': -2538}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011011; Y = 8'b10100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1283,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2538
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b10101110; // Expected: {'Z': -8446}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b10101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1284,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8446
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000110; Y = 8'b10011101; // Expected: {'Z': 5742}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000110; Y = 8'b10011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1285,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5742
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b01101100; // Expected: {'Z': 1404}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b01101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1286,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1404
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010010; Y = 8'b01000000; // Expected: {'Z': 5248}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010010; Y = 8'b01000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1287,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101011; Y = 8'b01011011; // Expected: {'Z': 3913}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101011; Y = 8'b01011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1288,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3913
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101000; Y = 8'b10000000; // Expected: {'Z': -5120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101000; Y = 8'b10000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1289,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b00111011; // Expected: {'Z': 1298}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b00111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1290,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1298
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b10110011; // Expected: {'Z': -1694}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b10110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1291,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1694
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100111; Y = 8'b11101110; // Expected: {'Z': 1602}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100111; Y = 8'b11101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1292,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1602
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010101; Y = 8'b00000010; // Expected: {'Z': 170}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010101; Y = 8'b00000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1293,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000111; Y = 8'b11011001; // Expected: {'Z': -2769}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000111; Y = 8'b11011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1294,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2769
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b01010100; // Expected: {'Z': 3276}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b01010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1295,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3276
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000000; Y = 8'b01011001; // Expected: {'Z': 5696}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000000; Y = 8'b01011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1296,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5696
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000000; Y = 8'b11010010; // Expected: {'Z': 5888}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000000; Y = 8'b11010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1297,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111101; Y = 8'b11011110; // Expected: {'Z': 2278}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111101; Y = 8'b11011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1298,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2278
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b00001000; // Expected: {'Z': 896}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b00001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1299,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b00011111; // Expected: {'Z': 899}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b00011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1300,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 899
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111110; Y = 8'b01010111; // Expected: {'Z': -5742}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111110; Y = 8'b01010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1301,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5742
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b11111010; // Expected: {'Z': -132}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b11111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1302,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b00011010; // Expected: {'Z': 1404}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b00011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1303,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1404
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b10101110; // Expected: {'Z': -3854}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b10101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1304,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3854
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111011; Y = 8'b00110001; // Expected: {'Z': -3381}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111011; Y = 8'b00110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1305,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3381
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010100; Y = 8'b01001000; // Expected: {'Z': -3168}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010100; Y = 8'b01001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1306,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000111; Y = 8'b10010000; // Expected: {'Z': -784}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000111; Y = 8'b10010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1307,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b00111100; // Expected: {'Z': 1260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b00111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1308,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101110; Y = 8'b11100011; // Expected: {'Z': -3190}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101110; Y = 8'b11100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1309,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b10110111; // Expected: {'Z': -7008}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b10110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1310,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b11011100; // Expected: {'Z': -1584}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b11011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1311,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1584
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000110; Y = 8'b11100111; // Expected: {'Z': 3050}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000110; Y = 8'b11100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1312,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100101; Y = 8'b01111110; // Expected: {'Z': 12726}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100101; Y = 8'b01111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1313,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 12726
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b11110010; // Expected: {'Z': -1722}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b11110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1314,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1722
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111001; Y = 8'b11011001; // Expected: {'Z': -2223}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111001; Y = 8'b11011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1315,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2223
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011011; Y = 8'b11011010; // Expected: {'Z': 1406}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011011; Y = 8'b11011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1316,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1406
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000111; Y = 8'b00100010; // Expected: {'Z': -4114}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000111; Y = 8'b00100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1317,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b11111011; // Expected: {'Z': -105}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b11111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1318,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011010; Y = 8'b01010010; // Expected: {'Z': -8364}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011010; Y = 8'b01010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1319,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010111; Y = 8'b01101011; // Expected: {'Z': -4387}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010111; Y = 8'b01101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1320,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4387
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101010; Y = 8'b00111001; // Expected: {'Z': -1254}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101010; Y = 8'b00111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1321,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110010; Y = 8'b10000000; // Expected: {'Z': 1792}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110010; Y = 8'b10000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1322,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000011; Y = 8'b10101111; // Expected: {'Z': -243}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000011; Y = 8'b10101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1323,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110011; Y = 8'b11110010; // Expected: {'Z': -1610}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110011; Y = 8'b11110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1324,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1610
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011110; Y = 8'b01011101; // Expected: {'Z': -3162}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011110; Y = 8'b01011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1325,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100101; Y = 8'b11000011; // Expected: {'Z': -2257}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100101; Y = 8'b11000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1326,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2257
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b11011000; // Expected: {'Z': 3360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b11011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1327,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001100; Y = 8'b10101011; // Expected: {'Z': 4420}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001100; Y = 8'b10101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1328,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111111; Y = 8'b11110011; // Expected: {'Z': -819}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111111; Y = 8'b11110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1329,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -819
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b00000101; // Expected: {'Z': 370}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b00000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1330,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 370
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b01001001; // Expected: {'Z': 2117}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b01001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1331,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110101; Y = 8'b00000101; // Expected: {'Z': 585}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110101; Y = 8'b00000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1332,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 585
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100010; Y = 8'b10100110; // Expected: {'Z': 8460}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100010; Y = 8'b10100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1333,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8460
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010011; Y = 8'b00001010; // Expected: {'Z': -450}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010011; Y = 8'b00001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1334,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111010; Y = 8'b10010110; // Expected: {'Z': 636}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111010; Y = 8'b10010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1335,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 636
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100110; Y = 8'b01111111; // Expected: {'Z': -11430}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100110; Y = 8'b01111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1336,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000110; Y = 8'b11011111; // Expected: {'Z': 4026}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000110; Y = 8'b11011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1337,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4026
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b11010101; // Expected: {'Z': 2408}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b11010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1338,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001011; Y = 8'b00000001; // Expected: {'Z': -53}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001011; Y = 8'b00000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1339,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b00101101; // Expected: {'Z': -1260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b00101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1340,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110110; Y = 8'b00010111; // Expected: {'Z': 2714}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110110; Y = 8'b00010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1341,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2714
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000011; Y = 8'b11011000; // Expected: {'Z': 2440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000011; Y = 8'b11011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1342,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b10100000; // Expected: {'Z': -2784}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b10100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1343,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101101; Y = 8'b01101001; // Expected: {'Z': -8715}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101101; Y = 8'b01101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1344,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8715
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010011; Y = 8'b00100100; // Expected: {'Z': 2988}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010011; Y = 8'b00100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1345,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2988
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b10101011; // Expected: {'Z': 5015}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b10101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1346,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5015
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110010; Y = 8'b01001010; // Expected: {'Z': 8436}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110010; Y = 8'b01001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1347,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8436
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000110; Y = 8'b01100010; // Expected: {'Z': -5684}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000110; Y = 8'b01100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1348,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5684
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100000; Y = 8'b11001001; // Expected: {'Z': -1760}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100000; Y = 8'b11001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1349,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110011; Y = 8'b10010001; // Expected: {'Z': -12765}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110011; Y = 8'b10010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1350,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12765
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000011; Y = 8'b00111111; // Expected: {'Z': 189}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000011; Y = 8'b00111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1351,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101000; Y = 8'b11010101; // Expected: {'Z': 3784}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101000; Y = 8'b11010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1352,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100110; Y = 8'b01001101; // Expected: {'Z': -6930}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100110; Y = 8'b01001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1353,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6930
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010111; Y = 8'b10100011; // Expected: {'Z': -8091}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010111; Y = 8'b10100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1354,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8091
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b00000001; // Expected: {'Z': 112}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b00000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1355,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b00011001; // Expected: {'Z': -1275}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b00011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1356,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1275
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001000; Y = 8'b10101111; // Expected: {'Z': 9720}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001000; Y = 8'b10101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1357,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b01101100; // Expected: {'Z': 10368}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b01101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1358,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101001; Y = 8'b00111110; // Expected: {'Z': 6510}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101001; Y = 8'b00111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1359,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6510
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000101; Y = 8'b11110111; // Expected: {'Z': -621}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000101; Y = 8'b11110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1360,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -621
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b11011110; // Expected: {'Z': -204}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b11011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1361,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101101; Y = 8'b11010101; // Expected: {'Z': 817}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101101; Y = 8'b11010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1362,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 817
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010100; Y = 8'b00011000; // Expected: {'Z': 2016}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010100; Y = 8'b00011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1363,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011001; Y = 8'b00111000; // Expected: {'Z': 4984}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011001; Y = 8'b00111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1364,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4984
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111100; Y = 8'b11011001; // Expected: {'Z': 156}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111100; Y = 8'b11011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1365,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100001; Y = 8'b11001101; // Expected: {'Z': -4947}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100001; Y = 8'b11001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1366,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4947
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110010; Y = 8'b10010111; // Expected: {'Z': 8190}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110010; Y = 8'b10010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1367,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b00100101; // Expected: {'Z': -3034}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b00100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1368,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3034
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110110; Y = 8'b00110001; // Expected: {'Z': -490}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110110; Y = 8'b00110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1369,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -490
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b11000000; // Expected: {'Z': 5376}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b11000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1370,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5376
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b01110000; // Expected: {'Z': 1680}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b01110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1371,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100010; Y = 8'b10111000; // Expected: {'Z': -2448}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100010; Y = 8'b10111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1372,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2448
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001101; Y = 8'b01011000; // Expected: {'Z': 6776}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001101; Y = 8'b01011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1373,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6776
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110101; Y = 8'b10001011; // Expected: {'Z': -6201}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110101; Y = 8'b10001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1374,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111111; Y = 8'b00011011; // Expected: {'Z': -1755}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111111; Y = 8'b00011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1375,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1755
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b01100101; // Expected: {'Z': 606}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b01100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1376,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 606
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001100; Y = 8'b01101000; // Expected: {'Z': -12064}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001100; Y = 8'b01101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1377,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12064
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101101; Y = 8'b00100111; // Expected: {'Z': 1755}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101101; Y = 8'b00100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1378,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1755
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000110; Y = 8'b01000010; // Expected: {'Z': -3828}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000110; Y = 8'b01000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1379,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110001; Y = 8'b00111010; // Expected: {'Z': 6554}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110001; Y = 8'b00111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1380,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6554
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111111; Y = 8'b01111110; // Expected: {'Z': -126}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111111; Y = 8'b01111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1381,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b10101110; // Expected: {'Z': -5002}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b10101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1382,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5002
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001001; Y = 8'b10101011; // Expected: {'Z': -6205}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001001; Y = 8'b10101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1383,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011010; Y = 8'b01001011; // Expected: {'Z': -7650}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011010; Y = 8'b01001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1384,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100000; Y = 8'b00011110; // Expected: {'Z': -960}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100000; Y = 8'b00011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1385,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001001; Y = 8'b00010001; // Expected: {'Z': -935}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001001; Y = 8'b00010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1386,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -935
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000101; Y = 8'b11101010; // Expected: {'Z': 2706}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000101; Y = 8'b11101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1387,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2706
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011000; Y = 8'b01101111; // Expected: {'Z': -11544}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011000; Y = 8'b01101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1388,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11544
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011011; Y = 8'b01001111; // Expected: {'Z': 7189}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011011; Y = 8'b01001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1389,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001110; Y = 8'b00011000; // Expected: {'Z': -1200}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001110; Y = 8'b00011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1390,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b00110100; // Expected: {'Z': 2444}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b00110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1391,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2444
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001000; Y = 8'b01110011; // Expected: {'Z': -13800}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001000; Y = 8'b01110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1392,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -13800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010111; Y = 8'b11110011; // Expected: {'Z': -299}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010111; Y = 8'b11110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1393,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -299
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010000; Y = 8'b00001100; // Expected: {'Z': -576}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010000; Y = 8'b00001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1394,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110101; Y = 8'b11111100; // Expected: {'Z': 44}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110101; Y = 8'b11111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1395,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100110; Y = 8'b11101011; // Expected: {'Z': -798}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100110; Y = 8'b11101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1396,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001111; Y = 8'b10111001; // Expected: {'Z': 8023}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001111; Y = 8'b10111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1397,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8023
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011001; Y = 8'b11101010; // Expected: {'Z': -1958}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011001; Y = 8'b11101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1398,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1958
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100101; Y = 8'b11111111; // Expected: {'Z': -37}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100101; Y = 8'b11111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1399,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110101; Y = 8'b00000100; // Expected: {'Z': 468}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110101; Y = 8'b00000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1400,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 468
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110100; Y = 8'b00100110; // Expected: {'Z': -2888}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110100; Y = 8'b00100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1401,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011011; Y = 8'b11101101; // Expected: {'Z': 1919}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011011; Y = 8'b11101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1402,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1919
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111011; Y = 8'b10100000; // Expected: {'Z': -5664}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111011; Y = 8'b10100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1403,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5664
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010100; Y = 8'b11101000; // Expected: {'Z': 2592}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010100; Y = 8'b11101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1404,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2592
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010110; Y = 8'b11011000; // Expected: {'Z': -3440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010110; Y = 8'b11011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1405,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b11101110; // Expected: {'Z': -1098}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b11101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1406,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1098
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b10110101; // Expected: {'Z': -1125}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b10110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1407,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b10100010; // Expected: {'Z': -3666}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b10100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1408,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3666
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001100; Y = 8'b10000100; // Expected: {'Z': -1488}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001100; Y = 8'b10000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1409,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101010; Y = 8'b00000010; // Expected: {'Z': -172}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101010; Y = 8'b00000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1410,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101010; Y = 8'b00110000; // Expected: {'Z': 5088}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101010; Y = 8'b00110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1411,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5088
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101111; Y = 8'b11110001; // Expected: {'Z': 1215}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101111; Y = 8'b11110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1412,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1215
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111101; Y = 8'b10110110; // Expected: {'Z': 4958}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111101; Y = 8'b10110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1413,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4958
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110011; Y = 8'b10011010; // Expected: {'Z': -11730}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110011; Y = 8'b10011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1414,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11730
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b00100101; // Expected: {'Z': 2516}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b00100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1415,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2516
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000001; Y = 8'b01001000; // Expected: {'Z': 4680}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000001; Y = 8'b01001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1416,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010010; Y = 8'b11110101; // Expected: {'Z': -198}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010010; Y = 8'b11110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1417,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010110; Y = 8'b01110110; // Expected: {'Z': 10148}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010110; Y = 8'b01110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1418,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000100; Y = 8'b01010100; // Expected: {'Z': -10416}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000100; Y = 8'b01010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1419,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111000; Y = 8'b01001101; // Expected: {'Z': 9240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111000; Y = 8'b01001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1420,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111011; Y = 8'b11100000; // Expected: {'Z': -1888}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111011; Y = 8'b11100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1421,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b01110111; // Expected: {'Z': 5236}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b01110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1422,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000000; Y = 8'b10001101; // Expected: {'Z': 7360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000000; Y = 8'b10001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1423,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011000; Y = 8'b01001011; // Expected: {'Z': -3000}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011000; Y = 8'b01001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1424,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010110; Y = 8'b00100010; // Expected: {'Z': -3604}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010110; Y = 8'b00100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1425,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3604
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000111; Y = 8'b10111011; // Expected: {'Z': -4899}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000111; Y = 8'b10111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1426,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4899
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b01010110; // Expected: {'Z': -4816}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b01010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1427,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000111; Y = 8'b10010100; // Expected: {'Z': 13068}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000111; Y = 8'b10010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1428,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 13068
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010000; Y = 8'b11000000; // Expected: {'Z': -5120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010000; Y = 8'b11000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1429,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100110; Y = 8'b00101010; // Expected: {'Z': -1092}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100110; Y = 8'b00101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1430,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1092
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011010; Y = 8'b11111110; // Expected: {'Z': -180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011010; Y = 8'b11111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1431,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100101; Y = 8'b01111100; // Expected: {'Z': 12524}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100101; Y = 8'b01111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1432,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 12524
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011010; Y = 8'b10101000; // Expected: {'Z': -7920}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011010; Y = 8'b10101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1433,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110001; Y = 8'b00000110; // Expected: {'Z': -474}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110001; Y = 8'b00000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1434,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -474
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011100; Y = 8'b00001001; // Expected: {'Z': -900}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011100; Y = 8'b00001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1435,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b11110100; // Expected: {'Z': -264}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b11110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1436,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101010; Y = 8'b10001011; // Expected: {'Z': -12402}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101010; Y = 8'b10001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1437,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12402
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010100; Y = 8'b00100001; // Expected: {'Z': -1452}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010100; Y = 8'b00100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1438,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1452
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100011; Y = 8'b00100111; // Expected: {'Z': 1365}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100011; Y = 8'b00100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1439,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1365
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110110; Y = 8'b10011011; // Expected: {'Z': 1010}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110110; Y = 8'b10011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1440,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1010
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101010; Y = 8'b00010100; // Expected: {'Z': 2120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101010; Y = 8'b00010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1441,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000010; Y = 8'b01001110; // Expected: {'Z': 5148}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000010; Y = 8'b01001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1442,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b11010101; // Expected: {'Z': -387}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b11010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1443,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -387
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010011; Y = 8'b00010110; // Expected: {'Z': 1826}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010011; Y = 8'b00010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1444,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1826
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111101; Y = 8'b00111010; // Expected: {'Z': 7250}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111101; Y = 8'b00111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1445,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000001; Y = 8'b10000000; // Expected: {'Z': -8320}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000001; Y = 8'b10000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1446,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000011; Y = 8'b01100010; // Expected: {'Z': 294}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000011; Y = 8'b01100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1447,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 294
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000000; Y = 8'b11111101; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000000; Y = 8'b11111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1448,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111001; Y = 8'b01111001; // Expected: {'Z': -847}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111001; Y = 8'b01111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1449,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -847
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000011; Y = 8'b01101100; // Expected: {'Z': -13500}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000011; Y = 8'b01101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1450,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -13500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111010; Y = 8'b01110010; // Expected: {'Z': 6612}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111010; Y = 8'b01110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1451,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100101; Y = 8'b00000010; // Expected: {'Z': -182}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100101; Y = 8'b00000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1452,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001110; Y = 8'b10000100; // Expected: {'Z': 6200}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001110; Y = 8'b10000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1453,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010101; Y = 8'b00000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010101; Y = 8'b00000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1454,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100011; Y = 8'b01111010; // Expected: {'Z': -11346}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100011; Y = 8'b01111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1455,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11346
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010100; Y = 8'b00001100; // Expected: {'Z': -528}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010100; Y = 8'b00001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1456,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b10110001; // Expected: {'Z': -1185}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b10110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1457,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011100; Y = 8'b01110111; // Expected: {'Z': 3332}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011100; Y = 8'b01110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1458,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3332
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b00111000; // Expected: {'Z': 4144}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b00111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1459,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101011; Y = 8'b01110110; // Expected: {'Z': 5074}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101011; Y = 8'b01110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1460,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5074
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100010; Y = 8'b10001110; // Expected: {'Z': -3876}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100010; Y = 8'b10001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1461,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3876
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110101; Y = 8'b00100000; // Expected: {'Z': 1696}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110101; Y = 8'b00100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1462,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1696
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101101; Y = 8'b01011011; // Expected: {'Z': 9919}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101101; Y = 8'b01011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1463,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9919
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001111; Y = 8'b01101001; // Expected: {'Z': -11865}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001111; Y = 8'b01101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1464,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11865
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011111; Y = 8'b10001111; // Expected: {'Z': 3729}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011111; Y = 8'b10001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1465,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3729
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110010; Y = 8'b11000001; // Expected: {'Z': -7182}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110010; Y = 8'b11000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1466,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100010; Y = 8'b00000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100010; Y = 8'b00000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1467,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000110; Y = 8'b01000001; // Expected: {'Z': -3770}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000110; Y = 8'b01000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1468,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3770
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b11100011; // Expected: {'Z': 3219}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b11100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1469,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3219
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011111; Y = 8'b01111101; // Expected: {'Z': -12125}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011111; Y = 8'b01111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1470,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b10000101; // Expected: {'Z': -246}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b10000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1471,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110111; Y = 8'b10011110; // Expected: {'Z': -11662}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110111; Y = 8'b10011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1472,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11662
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000110; Y = 8'b01011101; // Expected: {'Z': 6510}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000110; Y = 8'b01011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1473,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6510
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010100; Y = 8'b00110000; // Expected: {'Z': 960}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010100; Y = 8'b00110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1474,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100110; Y = 8'b10110010; // Expected: {'Z': 7020}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100110; Y = 8'b10110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1475,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7020
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011011; Y = 8'b00010100; // Expected: {'Z': -740}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011011; Y = 8'b00010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1476,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -740
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101010; Y = 8'b11000101; // Expected: {'Z': -6254}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101010; Y = 8'b11000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1477,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110100; Y = 8'b01111011; // Expected: {'Z': -9348}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110100; Y = 8'b01111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1478,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9348
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000001; Y = 8'b00000110; // Expected: {'Z': 390}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000001; Y = 8'b00000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1479,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 390
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011001; Y = 8'b11100110; // Expected: {'Z': 2678}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011001; Y = 8'b11100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1480,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2678
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111001; Y = 8'b10001101; // Expected: {'Z': -13915}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111001; Y = 8'b10001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1481,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -13915
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011001; Y = 8'b11000001; // Expected: {'Z': -1575}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011001; Y = 8'b11000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1482,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1575
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101100; Y = 8'b01001111; // Expected: {'Z': -1580}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101100; Y = 8'b01001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1483,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000000; Y = 8'b11111000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000000; Y = 8'b11111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1484,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110001; Y = 8'b10011110; // Expected: {'Z': 7742}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110001; Y = 8'b10011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1485,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7742
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100001; Y = 8'b01000011; // Expected: {'Z': -2077}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100001; Y = 8'b01000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1486,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2077
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010010; Y = 8'b01010001; // Expected: {'Z': -3726}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010010; Y = 8'b01010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1487,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3726
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010111; Y = 8'b00111001; // Expected: {'Z': 4959}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010111; Y = 8'b00111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1488,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4959
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011010; Y = 8'b11100001; // Expected: {'Z': -2790}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011010; Y = 8'b11100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1489,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2790
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b01101110; // Expected: {'Z': 3960}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b01101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1490,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b01001000; // Expected: {'Z': 2592}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b01001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1491,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2592
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b01010110; // Expected: {'Z': -4386}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b01010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1492,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4386
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110100; Y = 8'b01001010; // Expected: {'Z': 8584}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110100; Y = 8'b01001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1493,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8584
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111010; Y = 8'b01111110; // Expected: {'Z': -756}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111010; Y = 8'b01111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1494,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010011; Y = 8'b01011011; // Expected: {'Z': -4095}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010011; Y = 8'b01011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1495,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4095
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010000; Y = 8'b11010100; // Expected: {'Z': 4928}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010000; Y = 8'b11010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1496,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4928
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000000; Y = 8'b01001011; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000000; Y = 8'b01001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1497,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011011; Y = 8'b01110110; // Expected: {'Z': 10738}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011011; Y = 8'b01110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1498,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10738
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111010; Y = 8'b00000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111010; Y = 8'b00000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1499,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010010; Y = 8'b10100011; // Expected: {'Z': 4278}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010010; Y = 8'b10100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1500,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4278
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001010; Y = 8'b10100010; // Expected: {'Z': -940}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001010; Y = 8'b10100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1501,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -940
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010100; Y = 8'b10010011; // Expected: {'Z': -9156}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010100; Y = 8'b10010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1502,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000010; Y = 8'b00111101; // Expected: {'Z': -3782}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000010; Y = 8'b00111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1503,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3782
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011111; Y = 8'b11111000; // Expected: {'Z': 776}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011111; Y = 8'b11111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1504,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 776
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b00111000; // Expected: {'Z': 2632}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b00111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1505,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2632
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011100; Y = 8'b01100111; // Expected: {'Z': 2884}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011100; Y = 8'b01100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1506,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2884
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b10000100; // Expected: {'Z': 7316}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b10000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1507,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7316
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b10111110; // Expected: {'Z': -8118}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b10111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1508,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111110; Y = 8'b10101001; // Expected: {'Z': 174}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111110; Y = 8'b10101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1509,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000010; Y = 8'b01010011; // Expected: {'Z': -5146}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000010; Y = 8'b01010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1510,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b00100101; // Expected: {'Z': 1628}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b00100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1511,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1628
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101000; Y = 8'b00111101; // Expected: {'Z': 2440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101000; Y = 8'b00111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1512,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110001; Y = 8'b10010011; // Expected: {'Z': 8611}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110001; Y = 8'b10010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1513,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8611
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110010; Y = 8'b01100010; // Expected: {'Z': -7644}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110010; Y = 8'b01100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1514,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7644
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001101; Y = 8'b11100111; // Expected: {'Z': 2875}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001101; Y = 8'b11100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1515,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2875
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111010; Y = 8'b01011001; // Expected: {'Z': -6230}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111010; Y = 8'b01011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1516,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000011; Y = 8'b10101000; // Expected: {'Z': 11000}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000011; Y = 8'b10101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1517,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001010; Y = 8'b11001111; // Expected: {'Z': -490}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001010; Y = 8'b11001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1518,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -490
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001011; Y = 8'b10110010; // Expected: {'Z': 9126}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001011; Y = 8'b10110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1519,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110011; Y = 8'b00001000; // Expected: {'Z': 920}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110011; Y = 8'b00001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1520,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b11000111; // Expected: {'Z': 3363}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b11000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1521,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3363
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001100; Y = 8'b10001000; // Expected: {'Z': -9120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001100; Y = 8'b10001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1522,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001000; Y = 8'b11010100; // Expected: {'Z': 5280}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001000; Y = 8'b11010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1523,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100001; Y = 8'b00101010; // Expected: {'Z': -1302}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100001; Y = 8'b00101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1524,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1302
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110010; Y = 8'b01000101; // Expected: {'Z': 3450}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110010; Y = 8'b01000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1525,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001110; Y = 8'b11001110; // Expected: {'Z': 5700}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001110; Y = 8'b11001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1526,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001111; Y = 8'b00100001; // Expected: {'Z': -1617}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001111; Y = 8'b00100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1527,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1617
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b10010111; // Expected: {'Z': -3780}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b10010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1528,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010010; Y = 8'b11111101; // Expected: {'Z': 138}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010010; Y = 8'b11111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1529,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100010; Y = 8'b01100001; // Expected: {'Z': 9506}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100010; Y = 8'b01100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1530,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9506
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011110; Y = 8'b10001001; // Expected: {'Z': 11662}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011110; Y = 8'b10001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1531,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11662
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011101; Y = 8'b11000110; // Expected: {'Z': 2030}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011101; Y = 8'b11000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1532,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2030
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010000; Y = 8'b00110111; // Expected: {'Z': 880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010000; Y = 8'b00110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1533,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011101; Y = 8'b01001000; // Expected: {'Z': -2520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011101; Y = 8'b01001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1534,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010100; Y = 8'b11101101; // Expected: {'Z': 2052}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010100; Y = 8'b11101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1535,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2052
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000111; Y = 8'b10100011; // Expected: {'Z': 5301}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000111; Y = 8'b10100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1536,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5301
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010110; Y = 8'b00011001; // Expected: {'Z': -1050}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010110; Y = 8'b00011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1537,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011110; Y = 8'b00010010; // Expected: {'Z': 540}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011110; Y = 8'b00010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1538,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011110; Y = 8'b00000010; // Expected: {'Z': 188}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011110; Y = 8'b00000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1539,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011111; Y = 8'b00000011; // Expected: {'Z': 285}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011111; Y = 8'b00000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1540,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 285
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101101; Y = 8'b11111101; // Expected: {'Z': 57}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101101; Y = 8'b11111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1541,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010100; Y = 8'b11111010; // Expected: {'Z': -120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010100; Y = 8'b11111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1542,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111101; Y = 8'b11011110; // Expected: {'Z': 102}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111101; Y = 8'b11011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1543,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010100; Y = 8'b01011001; // Expected: {'Z': 1780}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010100; Y = 8'b01011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1544,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111100; Y = 8'b11110100; // Expected: {'Z': 48}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111100; Y = 8'b11110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1545,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b10000111; // Expected: {'Z': -4356}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b10000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1546,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4356
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010101; Y = 8'b01001100; // Expected: {'Z': -8132}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010101; Y = 8'b01001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1547,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100101; Y = 8'b10111100; // Expected: {'Z': -2516}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100101; Y = 8'b10111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1548,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2516
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111000; Y = 8'b11011000; // Expected: {'Z': -4800}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111000; Y = 8'b11011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1549,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100100; Y = 8'b01100001; // Expected: {'Z': -8924}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100100; Y = 8'b01100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1550,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8924
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001011; Y = 8'b10011000; // Expected: {'Z': 5512}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001011; Y = 8'b10011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1551,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5512
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101101; Y = 8'b10010101; // Expected: {'Z': 2033}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101101; Y = 8'b10010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1552,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2033
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b00100101; // Expected: {'Z': 4551}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b00100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1553,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4551
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000010; Y = 8'b10101010; // Expected: {'Z': 5332}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000010; Y = 8'b10101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1554,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5332
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000010; Y = 8'b10011100; // Expected: {'Z': 12600}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000010; Y = 8'b10011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1555,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 12600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101001; Y = 8'b00110000; // Expected: {'Z': 5040}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101001; Y = 8'b00110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1556,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111001; Y = 8'b10010100; // Expected: {'Z': -13068}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111001; Y = 8'b10010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1557,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -13068
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110001; Y = 8'b10111111; // Expected: {'Z': -7345}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110001; Y = 8'b10111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1558,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7345
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100011; Y = 8'b10011000; // Expected: {'Z': -10296}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100011; Y = 8'b10011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1559,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b10110100; // Expected: {'Z': -5472}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b10110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1560,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5472
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111110; Y = 8'b10101111; // Expected: {'Z': -5022}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111110; Y = 8'b10101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1561,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5022
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101111; Y = 8'b10111101; // Expected: {'Z': 5427}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101111; Y = 8'b10111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1562,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5427
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011100; Y = 8'b01011110; // Expected: {'Z': -3384}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011100; Y = 8'b01011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1563,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3384
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100000; Y = 8'b00010110; // Expected: {'Z': -2112}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100000; Y = 8'b00010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1564,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b01010001; // Expected: {'Z': -8991}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b01010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1565,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8991
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010100; Y = 8'b11000010; // Expected: {'Z': -5208}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010100; Y = 8'b11000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1566,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000011; Y = 8'b00000110; // Expected: {'Z': -366}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000011; Y = 8'b00000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1567,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -366
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101010; Y = 8'b10100110; // Expected: {'Z': -9540}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101010; Y = 8'b10100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1568,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110101; Y = 8'b01110101; // Expected: {'Z': -1287}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110101; Y = 8'b01110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1569,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1287
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b10011011; // Expected: {'Z': -4747}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b10011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1570,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4747
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b10100010; // Expected: {'Z': 8178}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b10100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1571,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111101; Y = 8'b00100110; // Expected: {'Z': 4750}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111101; Y = 8'b00100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1572,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001001; Y = 8'b10110000; // Expected: {'Z': 4400}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001001; Y = 8'b10110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1573,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101100; Y = 8'b10110110; // Expected: {'Z': 1480}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101100; Y = 8'b10110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1574,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111001; Y = 8'b11101011; // Expected: {'Z': -2541}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111001; Y = 8'b11101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1575,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2541
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b00111101; // Expected: {'Z': -5002}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b00111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1576,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5002
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110100; Y = 8'b11111101; // Expected: {'Z': 228}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110100; Y = 8'b11111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1577,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b10010001; // Expected: {'Z': -4884}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b10010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1578,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4884
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000001; Y = 8'b10011100; // Expected: {'Z': 6300}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000001; Y = 8'b10011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1579,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010101; Y = 8'b11000010; // Expected: {'Z': -5270}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010101; Y = 8'b11000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1580,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5270
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111101; Y = 8'b00011001; // Expected: {'Z': -75}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111101; Y = 8'b00011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1581,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110101; Y = 8'b00111111; // Expected: {'Z': -4725}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110101; Y = 8'b00111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1582,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4725
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010111; Y = 8'b01101110; // Expected: {'Z': -4510}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010111; Y = 8'b01101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1583,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4510
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010011; Y = 8'b11001001; // Expected: {'Z': -4565}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010011; Y = 8'b11001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1584,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4565
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011110; Y = 8'b10100001; // Expected: {'Z': -2850}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011110; Y = 8'b10100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1585,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2850
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010101; Y = 8'b00110111; // Expected: {'Z': -2365}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010101; Y = 8'b00110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1586,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2365
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111000; Y = 8'b11011111; // Expected: {'Z': -1848}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111000; Y = 8'b11011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1587,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010101; Y = 8'b00000001; // Expected: {'Z': -43}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010101; Y = 8'b00000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1588,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001000; Y = 8'b00000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001000; Y = 8'b00000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1589,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111010; Y = 8'b11000000; // Expected: {'Z': -7808}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111010; Y = 8'b11000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1590,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111011; Y = 8'b10111100; // Expected: {'Z': 4692}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111011; Y = 8'b10111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1591,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4692
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010001; Y = 8'b10101111; // Expected: {'Z': 3807}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010001; Y = 8'b10101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1592,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3807
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010010; Y = 8'b00110100; // Expected: {'Z': 4264}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010010; Y = 8'b00110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1593,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000010; Y = 8'b10000000; // Expected: {'Z': 16128}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000010; Y = 8'b10000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1594,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 16128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011101; Y = 8'b11110011; // Expected: {'Z': 455}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011101; Y = 8'b11110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1595,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 455
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110000; Y = 8'b00111011; // Expected: {'Z': -4720}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110000; Y = 8'b00111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1596,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110001; Y = 8'b10010101; // Expected: {'Z': 1605}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110001; Y = 8'b10010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1597,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1605
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010100; Y = 8'b11010001; // Expected: {'Z': -3948}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010100; Y = 8'b11010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1598,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3948
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110011; Y = 8'b01010001; // Expected: {'Z': 9315}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110011; Y = 8'b01010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1599,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9315
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110101; Y = 8'b00100010; // Expected: {'Z': -2550}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110101; Y = 8'b00100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1600,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011000; Y = 8'b00001110; // Expected: {'Z': -560}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011000; Y = 8'b00001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1601,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011001; Y = 8'b11101110; // Expected: {'Z': 702}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011001; Y = 8'b11101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1602,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 702
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b11000111; // Expected: {'Z': -342}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b11000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1603,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -342
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110010; Y = 8'b10111111; // Expected: {'Z': 5070}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110010; Y = 8'b10111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1604,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5070
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b00000001; // Expected: {'Z': 36}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b00000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1605,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011001; Y = 8'b10101110; // Expected: {'Z': -2050}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011001; Y = 8'b10101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1606,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110100; Y = 8'b00111001; // Expected: {'Z': 6612}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110100; Y = 8'b00111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1607,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110010; Y = 8'b00111011; // Expected: {'Z': -4602}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110010; Y = 8'b00111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1608,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4602
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101111; Y = 8'b00101011; // Expected: {'Z': -3483}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101111; Y = 8'b00101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1609,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3483
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001000; Y = 8'b01111001; // Expected: {'Z': 968}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001000; Y = 8'b01111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1610,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 968
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110011; Y = 8'b11010111; // Expected: {'Z': -4715}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110011; Y = 8'b11010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1611,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4715
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b10000111; // Expected: {'Z': -726}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b10000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1612,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -726
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010000; Y = 8'b11001110; // Expected: {'Z': -4000}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010000; Y = 8'b11001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1613,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100000; Y = 8'b01010010; // Expected: {'Z': -2624}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100000; Y = 8'b01010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1614,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111110; Y = 8'b00101101; // Expected: {'Z': -2970}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111110; Y = 8'b00101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1615,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2970
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000100; Y = 8'b00110101; // Expected: {'Z': 212}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000100; Y = 8'b00110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1616,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010110; Y = 8'b01100110; // Expected: {'Z': -4284}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010110; Y = 8'b01100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1617,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4284
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100110; Y = 8'b00100001; // Expected: {'Z': 3366}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100110; Y = 8'b00100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1618,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3366
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010010; Y = 8'b01110000; // Expected: {'Z': -12320}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010010; Y = 8'b01110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1619,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b11111011; // Expected: {'Z': 140}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b11111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1620,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b01110011; // Expected: {'Z': 5060}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b01110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1621,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010101; Y = 8'b01110010; // Expected: {'Z': -4902}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010101; Y = 8'b01110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1622,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4902
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110001; Y = 8'b11011010; // Expected: {'Z': 570}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110001; Y = 8'b11011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1623,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 570
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110100; Y = 8'b00101111; // Expected: {'Z': 5452}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110100; Y = 8'b00101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1624,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5452
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001010; Y = 8'b01001101; // Expected: {'Z': -9086}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001010; Y = 8'b01001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1625,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9086
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001110; Y = 8'b01110010; // Expected: {'Z': -5700}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001110; Y = 8'b01110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1626,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101010; Y = 8'b11101100; // Expected: {'Z': 1720}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101010; Y = 8'b11101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1627,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011011; Y = 8'b00011110; // Expected: {'Z': 810}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011011; Y = 8'b00011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1628,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 810
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100110; Y = 8'b10011010; // Expected: {'Z': 2652}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100110; Y = 8'b10011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1629,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2652
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b11001100; // Expected: {'Z': -3172}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b11001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1630,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100110; Y = 8'b01000011; // Expected: {'Z': -6030}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100110; Y = 8'b01000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1631,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6030
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110110; Y = 8'b10100011; // Expected: {'Z': 6882}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110110; Y = 8'b10100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1632,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6882
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100001; Y = 8'b11011111; // Expected: {'Z': 3135}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100001; Y = 8'b11011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1633,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b00011010; // Expected: {'Z': 1144}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b00011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1634,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b10100000; // Expected: {'Z': -6528}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b10100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1635,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101001; Y = 8'b10001100; // Expected: {'Z': -12180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101001; Y = 8'b10001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1636,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b01010111; // Expected: {'Z': -2436}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b01010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1637,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2436
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101110; Y = 8'b01111011; // Expected: {'Z': 13530}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101110; Y = 8'b01111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1638,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 13530
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111001; Y = 8'b11111110; // Expected: {'Z': -114}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111001; Y = 8'b11111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1639,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011010; Y = 8'b00010110; // Expected: {'Z': 572}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011010; Y = 8'b00010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1640,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 572
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111010; Y = 8'b10110101; // Expected: {'Z': -9150}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111010; Y = 8'b10110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1641,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000000; Y = 8'b01101110; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000000; Y = 8'b01101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1642,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010000; Y = 8'b11010110; // Expected: {'Z': 4704}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010000; Y = 8'b11010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1643,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4704
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011100; Y = 8'b00010100; // Expected: {'Z': 560}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011100; Y = 8'b00010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1644,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110111; Y = 8'b01101110; // Expected: {'Z': -990}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110111; Y = 8'b01101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1645,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -990
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001100; Y = 8'b00010100; // Expected: {'Z': 240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001100; Y = 8'b00010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1646,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001000; Y = 8'b11101011; // Expected: {'Z': -168}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001000; Y = 8'b11101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1647,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111000; Y = 8'b01100001; // Expected: {'Z': 11640}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111000; Y = 8'b01100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1648,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011100; Y = 8'b11110110; // Expected: {'Z': 1000}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011100; Y = 8'b11110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1649,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110111; Y = 8'b10110111; // Expected: {'Z': 5329}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110111; Y = 8'b10110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1650,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5329
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011111; Y = 8'b00011000; // Expected: {'Z': -2328}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011111; Y = 8'b00011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1651,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2328
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010011; Y = 8'b01101010; // Expected: {'Z': -11554}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010011; Y = 8'b01101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1652,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11554
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011100; Y = 8'b10001000; // Expected: {'Z': 4320}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011100; Y = 8'b10001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1653,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001100; Y = 8'b11010100; // Expected: {'Z': -528}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001100; Y = 8'b11010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1654,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010111; Y = 8'b10101101; // Expected: {'Z': 8715}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010111; Y = 8'b10101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1655,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8715
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111011; Y = 8'b10000111; // Expected: {'Z': -7139}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111011; Y = 8'b10000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1656,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7139
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b01100001; // Expected: {'Z': 9312}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b01100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1657,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9312
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001011; Y = 8'b00111011; // Expected: {'Z': -3127}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001011; Y = 8'b00111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1658,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3127
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010000; Y = 8'b00000001; // Expected: {'Z': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010000; Y = 8'b00000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1659,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110111; Y = 8'b11000101; // Expected: {'Z': 4307}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110111; Y = 8'b11000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1660,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4307
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100010; Y = 8'b01000100; // Expected: {'Z': -2040}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100010; Y = 8'b01000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1661,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b00111101; // Expected: {'Z': 3294}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b00111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1662,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3294
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110011; Y = 8'b00101111; // Expected: {'Z': -3619}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110011; Y = 8'b00101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1663,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3619
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110010; Y = 8'b00001111; // Expected: {'Z': -210}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110010; Y = 8'b00001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1664,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101100; Y = 8'b01110111; // Expected: {'Z': 12852}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101100; Y = 8'b01110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1665,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 12852
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111011; Y = 8'b01001111; // Expected: {'Z': -5451}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111011; Y = 8'b01001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1666,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5451
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001010; Y = 8'b01101011; // Expected: {'Z': -5778}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001010; Y = 8'b01101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1667,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5778
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000000; Y = 8'b10101010; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000000; Y = 8'b10101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1668,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110110; Y = 8'b01001100; // Expected: {'Z': -760}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110110; Y = 8'b01001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1669,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110111; Y = 8'b10001001; // Expected: {'Z': 8687}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110111; Y = 8'b10001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1670,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8687
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111011; Y = 8'b10100111; // Expected: {'Z': 6141}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111011; Y = 8'b10100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1671,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b10111010; // Expected: {'Z': -3080}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b10111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1672,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000001; Y = 8'b00100000; // Expected: {'Z': -4064}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000001; Y = 8'b00100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1673,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4064
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101100; Y = 8'b10100101; // Expected: {'Z': -9828}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101100; Y = 8'b10100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1674,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111011; Y = 8'b10010110; // Expected: {'Z': 530}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111011; Y = 8'b10010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1675,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 530
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010010; Y = 8'b00011010; // Expected: {'Z': 468}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010010; Y = 8'b00011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1676,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 468
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b00010101; // Expected: {'Z': 2163}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b00010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1677,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2163
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000100; Y = 8'b11100111; // Expected: {'Z': 1500}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000100; Y = 8'b11100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1678,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000001; Y = 8'b00111111; // Expected: {'Z': 4095}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000001; Y = 8'b00111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1679,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4095
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010100; Y = 8'b01000110; // Expected: {'Z': 1400}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010100; Y = 8'b01000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1680,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010101; Y = 8'b10101001; // Expected: {'Z': -7395}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010101; Y = 8'b10101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1681,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7395
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111111; Y = 8'b11100110; // Expected: {'Z': -3302}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111111; Y = 8'b11100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1682,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3302
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111010; Y = 8'b00100110; // Expected: {'Z': -228}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111010; Y = 8'b00100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1683,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010101; Y = 8'b01011011; // Expected: {'Z': -9737}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010101; Y = 8'b01011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1684,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9737
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100011; Y = 8'b01001100; // Expected: {'Z': -7068}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100011; Y = 8'b01001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1685,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7068
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110010; Y = 8'b01000000; // Expected: {'Z': -4992}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110010; Y = 8'b01000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1686,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4992
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001010; Y = 8'b10000100; // Expected: {'Z': -1240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001010; Y = 8'b10000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1687,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111011; Y = 8'b01111000; // Expected: {'Z': -8280}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111011; Y = 8'b01111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1688,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100110; Y = 8'b11001011; // Expected: {'Z': 4770}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100110; Y = 8'b11001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1689,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4770
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111111; Y = 8'b00010001; // Expected: {'Z': 2159}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111111; Y = 8'b00010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1690,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b01100000; // Expected: {'Z': 11808}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b01100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1691,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110000; Y = 8'b00010011; // Expected: {'Z': -304}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110000; Y = 8'b00010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1692,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -304
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001000; Y = 8'b11101100; // Expected: {'Z': -160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001000; Y = 8'b11101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1693,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101011; Y = 8'b11001000; // Expected: {'Z': -5992}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101011; Y = 8'b11001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1694,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5992
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b01110110; // Expected: {'Z': 5192}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b01110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1695,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101011; Y = 8'b10000000; // Expected: {'Z': 2688}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101011; Y = 8'b10000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1696,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2688
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b01000011; // Expected: {'Z': -4556}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b01000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1697,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4556
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011010; Y = 8'b10101010; // Expected: {'Z': -2236}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011010; Y = 8'b10101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1698,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011100; Y = 8'b01110011; // Expected: {'Z': -11500}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011100; Y = 8'b01110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1699,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011111; Y = 8'b00101110; // Expected: {'Z': -4462}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011111; Y = 8'b00101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1700,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000000; Y = 8'b11010011; // Expected: {'Z': -2880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000000; Y = 8'b11010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1701,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010001; Y = 8'b10100000; // Expected: {'Z': -1632}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010001; Y = 8'b10100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1702,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1632
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101110; Y = 8'b01010101; // Expected: {'Z': 9350}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101110; Y = 8'b01010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1703,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110101; Y = 8'b01011010; // Expected: {'Z': 10530}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110101; Y = 8'b01011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1704,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10530
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001101; Y = 8'b10000111; // Expected: {'Z': 13915}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001101; Y = 8'b10000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1705,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 13915
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111010; Y = 8'b01110001; // Expected: {'Z': 13786}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111010; Y = 8'b01110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1706,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 13786
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110110; Y = 8'b10000010; // Expected: {'Z': -14868}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110110; Y = 8'b10000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1707,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -14868
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011010; Y = 8'b11010011; // Expected: {'Z': -4050}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011010; Y = 8'b11010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1708,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b10000000; // Expected: {'Z': -12288}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b10000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1709,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001010; Y = 8'b00100010; // Expected: {'Z': 340}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001010; Y = 8'b00100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1710,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b11111111; // Expected: {'Z': -123}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b11111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1711,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -123
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011101; Y = 8'b10100100; // Expected: {'Z': -8556}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011101; Y = 8'b10100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1712,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8556
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b01101111; // Expected: {'Z': -7548}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b01101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1713,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7548
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000000; Y = 8'b10100000; // Expected: {'Z': 12288}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000000; Y = 8'b10100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1714,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 12288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111110; Y = 8'b10110010; // Expected: {'Z': -9828}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111110; Y = 8'b10110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1715,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110111; Y = 8'b01111011; // Expected: {'Z': 14637}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110111; Y = 8'b01111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1716,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 14637
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101001; Y = 8'b11001000; // Expected: {'Z': 1288}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101001; Y = 8'b11001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1717,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000101; Y = 8'b01111001; // Expected: {'Z': 605}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000101; Y = 8'b01111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1718,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 605
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010101; Y = 8'b10101100; // Expected: {'Z': 8988}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010101; Y = 8'b10101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1719,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8988
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101111; Y = 8'b01000001; // Expected: {'Z': 7215}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101111; Y = 8'b01000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1720,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7215
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001100; Y = 8'b01000100; // Expected: {'Z': -7888}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001100; Y = 8'b01000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1721,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110001; Y = 8'b01011011; // Expected: {'Z': -7189}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110001; Y = 8'b01011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1722,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100001; Y = 8'b01101011; // Expected: {'Z': 10379}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100001; Y = 8'b01101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1723,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10379
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000010; Y = 8'b01011110; // Expected: {'Z': 6204}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000010; Y = 8'b01011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1724,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000001; Y = 8'b00111010; // Expected: {'Z': 3770}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000001; Y = 8'b00111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1725,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3770
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010100; Y = 8'b10110010; // Expected: {'Z': 3432}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010100; Y = 8'b10110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1726,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000011; Y = 8'b11001000; // Expected: {'Z': 7000}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000011; Y = 8'b11001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1727,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000011; Y = 8'b10111110; // Expected: {'Z': -198}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000011; Y = 8'b10111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1728,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111011; Y = 8'b10111111; // Expected: {'Z': 325}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111011; Y = 8'b10111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1729,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 325
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110010; Y = 8'b10001001; // Expected: {'Z': 9282}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110010; Y = 8'b10001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1730,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9282
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100110; Y = 8'b01001001; // Expected: {'Z': -1898}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100110; Y = 8'b01001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1731,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1898
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101011; Y = 8'b00100011; // Expected: {'Z': 1505}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101011; Y = 8'b00100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1732,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1505
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000011; Y = 8'b01010000; // Expected: {'Z': -10000}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000011; Y = 8'b01010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1733,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011100; Y = 8'b01010111; // Expected: {'Z': -8700}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011100; Y = 8'b01010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1734,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000011; Y = 8'b00010111; // Expected: {'Z': 1541}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000011; Y = 8'b00010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1735,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1541
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111011; Y = 8'b10110001; // Expected: {'Z': 395}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111011; Y = 8'b10110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1736,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 395
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101011; Y = 8'b10110111; // Expected: {'Z': 6205}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101011; Y = 8'b10110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1737,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001111; Y = 8'b11111011; // Expected: {'Z': 245}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001111; Y = 8'b11111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1738,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b00111111; // Expected: {'Z': 378}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b00111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1739,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 378
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001100; Y = 8'b11001100; // Expected: {'Z': 6032}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001100; Y = 8'b11001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1740,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6032
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011101; Y = 8'b01001111; // Expected: {'Z': -7821}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011101; Y = 8'b01001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1741,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7821
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011100; Y = 8'b00000101; // Expected: {'Z': 460}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011100; Y = 8'b00000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1742,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 460
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b01111010; // Expected: {'Z': 7442}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b01111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1743,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7442
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101100; Y = 8'b01010101; // Expected: {'Z': -1700}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101100; Y = 8'b01010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1744,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100010; Y = 8'b00001111; // Expected: {'Z': -1410}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100010; Y = 8'b00001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1745,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1410
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001110; Y = 8'b10101100; // Expected: {'Z': -6552}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001110; Y = 8'b10101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1746,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b00101110; // Expected: {'Z': -3772}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b00101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1747,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3772
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000111; Y = 8'b11111001; // Expected: {'Z': -497}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000111; Y = 8'b11111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1748,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -497
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b11101010; // Expected: {'Z': 616}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b11101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1749,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 616
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111110; Y = 8'b01010011; // Expected: {'Z': -166}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111110; Y = 8'b01010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1750,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101111; Y = 8'b10010100; // Expected: {'Z': 1836}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101111; Y = 8'b10010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1751,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1836
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100010; Y = 8'b01101011; // Expected: {'Z': 10486}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100010; Y = 8'b01101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1752,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10486
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000111; Y = 8'b11101100; // Expected: {'Z': 2420}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000111; Y = 8'b11101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1753,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101010; Y = 8'b10100011; // Expected: {'Z': -9858}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101010; Y = 8'b10100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1754,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9858
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001100; Y = 8'b11000111; // Expected: {'Z': 6612}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001100; Y = 8'b11000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1755,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b11000000; // Expected: {'Z': 1792}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b11000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1756,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101010; Y = 8'b01111100; // Expected: {'Z': -2728}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101010; Y = 8'b01111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1757,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110001; Y = 8'b10001011; // Expected: {'Z': -13221}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110001; Y = 8'b10001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1758,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -13221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001100; Y = 8'b11011101; // Expected: {'Z': 1820}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001100; Y = 8'b11011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1759,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101000; Y = 8'b01110100; // Expected: {'Z': 12064}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101000; Y = 8'b01110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1760,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 12064
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001111; Y = 8'b10110110; // Expected: {'Z': 8362}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001111; Y = 8'b10110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1761,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8362
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011001; Y = 8'b10010110; // Expected: {'Z': 10918}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011001; Y = 8'b10010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1762,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10918
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011101; Y = 8'b00100011; // Expected: {'Z': -3465}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011101; Y = 8'b00100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1763,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3465
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001111; Y = 8'b10010101; // Expected: {'Z': 12091}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001111; Y = 8'b10010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1764,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 12091
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111111; Y = 8'b11111100; // Expected: {'Z': 260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111111; Y = 8'b11111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1765,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011111; Y = 8'b11000001; // Expected: {'Z': -5985}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011111; Y = 8'b11000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1766,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5985
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010010; Y = 8'b11110000; // Expected: {'Z': -288}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010010; Y = 8'b11110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1767,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101010; Y = 8'b10011010; // Expected: {'Z': 2244}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101010; Y = 8'b10011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1768,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000101; Y = 8'b11101110; // Expected: {'Z': -90}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000101; Y = 8'b11101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1769,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001111; Y = 8'b11100101; // Expected: {'Z': -2133}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001111; Y = 8'b11100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1770,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2133
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000100; Y = 8'b11100111; // Expected: {'Z': 3100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000100; Y = 8'b11100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1771,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000000; Y = 8'b00000011; // Expected: {'Z': -192}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000000; Y = 8'b00000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1772,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110101; Y = 8'b00100101; // Expected: {'Z': -407}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110101; Y = 8'b00100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1773,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -407
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101001; Y = 8'b01001100; // Expected: {'Z': -1748}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101001; Y = 8'b01001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1774,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1748
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011011; Y = 8'b10001101; // Expected: {'Z': 4255}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011011; Y = 8'b10001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1775,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110010; Y = 8'b11011100; // Expected: {'Z': 504}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110010; Y = 8'b11011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1776,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101100; Y = 8'b10101001; // Expected: {'Z': -9396}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101100; Y = 8'b10101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1777,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9396
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110101; Y = 8'b01101000; // Expected: {'Z': -7800}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110101; Y = 8'b01101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1778,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b10010001; // Expected: {'Z': 9324}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b10010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1779,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9324
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100000; Y = 8'b10110001; // Expected: {'Z': -2528}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100000; Y = 8'b10110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1780,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110110; Y = 8'b11011001; // Expected: {'Z': 390}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110110; Y = 8'b11011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1781,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 390
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b01111010; // Expected: {'Z': 9028}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b01111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1782,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9028
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100101; Y = 8'b11110101; // Expected: {'Z': 297}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100101; Y = 8'b11110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1783,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 297
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000000; Y = 8'b10110000; // Expected: {'Z': 5120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000000; Y = 8'b10110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1784,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000011; Y = 8'b10111000; // Expected: {'Z': -216}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000011; Y = 8'b10111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1785,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010000; Y = 8'b00101011; // Expected: {'Z': 3440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010000; Y = 8'b00101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1786,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011101; Y = 8'b01110101; // Expected: {'Z': 10881}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011101; Y = 8'b01110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1787,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10881
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010000; Y = 8'b10011011; // Expected: {'Z': -1616}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010000; Y = 8'b10011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1788,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1616
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010101; Y = 8'b01101111; // Expected: {'Z': 9435}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010101; Y = 8'b01101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1789,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9435
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010001; Y = 8'b01101010; // Expected: {'Z': 8586}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010001; Y = 8'b01101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1790,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8586
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000101; Y = 8'b10101111; // Expected: {'Z': -405}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000101; Y = 8'b10101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1791,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -405
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000011; Y = 8'b10010001; // Expected: {'Z': -7437}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000011; Y = 8'b10010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1792,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7437
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111111; Y = 8'b01010010; // Expected: {'Z': -5330}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111111; Y = 8'b01010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1793,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5330
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110110; Y = 8'b10100101; // Expected: {'Z': -10738}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110110; Y = 8'b10100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1794,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10738
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001000; Y = 8'b01110111; // Expected: {'Z': -14280}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001000; Y = 8'b01110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1795,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -14280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010000; Y = 8'b00101010; // Expected: {'Z': -2016}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010000; Y = 8'b00101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1796,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000111; Y = 8'b11011001; // Expected: {'Z': -273}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000111; Y = 8'b11011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1797,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -273
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010101; Y = 8'b10000001; // Expected: {'Z': 5461}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010101; Y = 8'b10000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1798,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5461
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101001; Y = 8'b01100010; // Expected: {'Z': -2254}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101001; Y = 8'b01100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1799,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000111; Y = 8'b00110111; // Expected: {'Z': 3905}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000111; Y = 8'b00110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1800,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3905
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010001; Y = 8'b01110111; // Expected: {'Z': 9639}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010001; Y = 8'b01110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1801,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9639
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000111; Y = 8'b10110110; // Expected: {'Z': 8954}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000111; Y = 8'b10110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1802,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8954
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010000; Y = 8'b10111101; // Expected: {'Z': -1072}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010000; Y = 8'b10111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1803,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1072
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b11111111; // Expected: {'Z': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b11111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1804,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011110; Y = 8'b00010000; // Expected: {'Z': 480}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011110; Y = 8'b00010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1805,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011010; Y = 8'b11011010; // Expected: {'Z': 1444}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011010; Y = 8'b11011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1806,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1444
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110010; Y = 8'b10010000; // Expected: {'Z': 1568}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110010; Y = 8'b10010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1807,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1568
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000011; Y = 8'b10111000; // Expected: {'Z': 9000}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000011; Y = 8'b10111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1808,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100101; Y = 8'b11101101; // Expected: {'Z': 513}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100101; Y = 8'b11101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1809,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 513
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011111; Y = 8'b10010101; // Expected: {'Z': 3531}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011111; Y = 8'b10010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1810,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3531
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110001; Y = 8'b00110000; // Expected: {'Z': 2352}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110001; Y = 8'b00110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1811,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001100; Y = 8'b00000001; // Expected: {'Z': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001100; Y = 8'b00000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1812,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111100; Y = 8'b11110110; // Expected: {'Z': 40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111100; Y = 8'b11110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1813,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011111; Y = 8'b01101100; // Expected: {'Z': -3564}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011111; Y = 8'b01101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1814,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3564
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101110; Y = 8'b11010101; // Expected: {'Z': -1978}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101110; Y = 8'b11010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1815,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1978
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b10000110; // Expected: {'Z': 10248}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b10000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1816,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b10011000; // Expected: {'Z': 7072}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b10011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1817,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7072
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010101; Y = 8'b10101110; // Expected: {'Z': -6970}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010101; Y = 8'b10101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1818,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6970
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100111; Y = 8'b10011010; // Expected: {'Z': 9078}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100111; Y = 8'b10011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1819,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9078
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b00111111; // Expected: {'Z': 7056}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b00111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1820,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7056
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011100; Y = 8'b01001100; // Expected: {'Z': -2736}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011100; Y = 8'b01001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1821,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000010; Y = 8'b10001110; // Expected: {'Z': 7068}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000010; Y = 8'b10001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1822,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7068
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010111; Y = 8'b00010011; // Expected: {'Z': 437}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010111; Y = 8'b00010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1823,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 437
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011001; Y = 8'b10010011; // Expected: {'Z': 11227}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011001; Y = 8'b10010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1824,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11227
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000010; Y = 8'b11110111; // Expected: {'Z': 1134}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000010; Y = 8'b11110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1825,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001011; Y = 8'b11011000; // Expected: {'Z': 4680}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001011; Y = 8'b11011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1826,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001110; Y = 8'b11011010; // Expected: {'Z': 1900}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001110; Y = 8'b11011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1827,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011001; Y = 8'b10101010; // Expected: {'Z': 3354}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011001; Y = 8'b10101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1828,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3354
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111001; Y = 8'b10000101; // Expected: {'Z': -7011}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111001; Y = 8'b10000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1829,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7011
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101010; Y = 8'b00100000; // Expected: {'Z': -2752}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101010; Y = 8'b00100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1830,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2752
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110000; Y = 8'b11110011; // Expected: {'Z': 1040}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110000; Y = 8'b11110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1831,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101101; Y = 8'b10110100; // Expected: {'Z': -8284}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101101; Y = 8'b10110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1832,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8284
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b10000110; // Expected: {'Z': -8296}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b10000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1833,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001011; Y = 8'b11001101; // Expected: {'Z': -3825}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001011; Y = 8'b11001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1834,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3825
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000100; Y = 8'b11110011; // Expected: {'Z': 780}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000100; Y = 8'b11110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1835,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011101; Y = 8'b10000111; // Expected: {'Z': -11253}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011101; Y = 8'b10000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1836,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b00010000; // Expected: {'Z': -816}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b00010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1837,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110000; Y = 8'b01111110; // Expected: {'Z': -2016}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110000; Y = 8'b01111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1838,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100011; Y = 8'b00000001; // Expected: {'Z': 99}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100011; Y = 8'b00000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1839,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110110; Y = 8'b10010111; // Expected: {'Z': -12390}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110110; Y = 8'b10010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1840,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12390
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000110; Y = 8'b11111011; // Expected: {'Z': -350}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000110; Y = 8'b11111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1841,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010100; Y = 8'b00101000; // Expected: {'Z': 800}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010100; Y = 8'b00101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1842,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100010; Y = 8'b10100101; // Expected: {'Z': 8554}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100010; Y = 8'b10100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1843,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8554
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010110; Y = 8'b00100111; // Expected: {'Z': -4134}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010110; Y = 8'b00100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1844,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001110; Y = 8'b11101000; // Expected: {'Z': -336}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001110; Y = 8'b11101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1845,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -336
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010000; Y = 8'b11001001; // Expected: {'Z': 6160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010000; Y = 8'b11001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1846,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010001; Y = 8'b11110111; // Expected: {'Z': 423}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010001; Y = 8'b11110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1847,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 423
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b01001110; // Expected: {'Z': 2262}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b01001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1848,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2262
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010001; Y = 8'b00100000; // Expected: {'Z': 2592}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010001; Y = 8'b00100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1849,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2592
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b01110001; // Expected: {'Z': -9492}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b01110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1850,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9492
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101101; Y = 8'b00011001; // Expected: {'Z': 1125}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101101; Y = 8'b00011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1851,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000011; Y = 8'b11111010; // Expected: {'Z': 750}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000011; Y = 8'b11111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1852,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110001; Y = 8'b01110111; // Expected: {'Z': -1785}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110001; Y = 8'b01110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1853,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1785
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111000; Y = 8'b10101100; // Expected: {'Z': 6048}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111000; Y = 8'b10101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1854,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6048
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100001; Y = 8'b01101111; // Expected: {'Z': 10767}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100001; Y = 8'b01101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1855,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10767
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011100; Y = 8'b11110110; // Expected: {'Z': -280}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011100; Y = 8'b11110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1856,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111010; Y = 8'b10000011; // Expected: {'Z': -15250}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111010; Y = 8'b10000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1857,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -15250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b10110001; // Expected: {'Z': -3081}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b10110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1858,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3081
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000000; Y = 8'b00100110; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000000; Y = 8'b00100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1859,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101000; Y = 8'b00111100; // Expected: {'Z': 6240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101000; Y = 8'b00111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1860,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100011; Y = 8'b00100001; // Expected: {'Z': 1155}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100011; Y = 8'b00100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1861,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101010; Y = 8'b00000101; // Expected: {'Z': -430}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101010; Y = 8'b00000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1862,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b10100011; // Expected: {'Z': -8928}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b10100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1863,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8928
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010010; Y = 8'b00101000; // Expected: {'Z': -1840}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010010; Y = 8'b00101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1864,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010001; Y = 8'b11111111; // Expected: {'Z': -81}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010001; Y = 8'b11111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1865,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b11000011; // Expected: {'Z': 6771}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b11000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1866,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6771
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001110; Y = 8'b01000111; // Expected: {'Z': -8094}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001110; Y = 8'b01000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1867,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8094
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100001; Y = 8'b10010101; // Expected: {'Z': -3531}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100001; Y = 8'b10010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1868,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3531
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101111; Y = 8'b10111111; // Expected: {'Z': 1105}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101111; Y = 8'b10111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1869,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b00001100; // Expected: {'Z': 156}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b00001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1870,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b11100001; // Expected: {'Z': -2728}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b11100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1871,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101101; Y = 8'b01110110; // Expected: {'Z': 12862}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101101; Y = 8'b01110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1872,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 12862
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b10010010; // Expected: {'Z': -7920}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b10010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1873,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101001; Y = 8'b11001011; // Expected: {'Z': -5565}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101001; Y = 8'b11001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1874,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5565
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b01011100; // Expected: {'Z': 8096}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b01011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1875,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8096
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b11011010; // Expected: {'Z': -2812}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b11011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1876,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2812
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b00001000; // Expected: {'Z': 168}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b00001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1877,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011000; Y = 8'b01100001; // Expected: {'Z': -10088}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011000; Y = 8'b01100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1878,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10088
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b00001011; // Expected: {'Z': -924}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b00001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1879,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -924
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b11010000; // Expected: {'Z': 2448}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b11010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1880,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2448
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000100; Y = 8'b01100001; // Expected: {'Z': -5820}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000100; Y = 8'b01100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1881,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000101; Y = 8'b00000101; // Expected: {'Z': 25}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000101; Y = 8'b00000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1882,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010110; Y = 8'b00000111; // Expected: {'Z': -294}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010110; Y = 8'b00000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1883,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -294
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101110; Y = 8'b01111011; // Expected: {'Z': -2214}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101110; Y = 8'b01111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1884,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000010; Y = 8'b01111111; // Expected: {'Z': 8382}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000010; Y = 8'b01111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1885,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8382
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011011; Y = 8'b00001101; // Expected: {'Z': -1313}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011011; Y = 8'b00001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1886,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1313
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111010; Y = 8'b11110101; // Expected: {'Z': -638}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111010; Y = 8'b11110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1887,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -638
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b10001000; // Expected: {'Z': -10560}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b10001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1888,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b00010011; // Expected: {'Z': -1558}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b00010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1889,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1558
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011010; Y = 8'b01011001; // Expected: {'Z': -3382}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011010; Y = 8'b01011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1890,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3382
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111110; Y = 8'b10101011; // Expected: {'Z': 170}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111110; Y = 8'b10101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1891,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b11110110; // Expected: {'Z': -680}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b11110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1892,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b10011110; // Expected: {'Z': -2156}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b10011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1893,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b01100100; // Expected: {'Z': -8200}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b01100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1894,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011111; Y = 8'b11100010; // Expected: {'Z': -2850}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011111; Y = 8'b11100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1895,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2850
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b00110100; // Expected: {'Z': 1508}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b00110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1896,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1508
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b00011111; // Expected: {'Z': 2728}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b00011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1897,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b00101110; // Expected: {'Z': 2806}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b00101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1898,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2806
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b10111110; // Expected: {'Z': -6336}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b10111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1899,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6336
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010010; Y = 8'b00011011; // Expected: {'Z': 2214}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010010; Y = 8'b00011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1900,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b01110010; // Expected: {'Z': 7752}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b01110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1901,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7752
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001011; Y = 8'b01000010; // Expected: {'Z': 726}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001011; Y = 8'b01000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1902,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 726
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101101; Y = 8'b01100011; // Expected: {'Z': 10791}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101101; Y = 8'b01100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1903,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10791
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000011; Y = 8'b00110101; // Expected: {'Z': -3233}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000011; Y = 8'b00110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1904,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3233
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100100; Y = 8'b10101010; // Expected: {'Z': -8600}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100100; Y = 8'b10101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1905,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011100; Y = 8'b11101001; // Expected: {'Z': 828}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011100; Y = 8'b11101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1906,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101010; Y = 8'b11101100; // Expected: {'Z': 440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101010; Y = 8'b11101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1907,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110100; Y = 8'b01010101; // Expected: {'Z': -6460}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110100; Y = 8'b01010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1908,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6460
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b10101000; // Expected: {'Z': 4488}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b10101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1909,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111101; Y = 8'b10000010; // Expected: {'Z': 378}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111101; Y = 8'b10000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1910,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 378
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010110; Y = 8'b10110001; // Expected: {'Z': 3318}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010110; Y = 8'b10110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1911,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3318
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110010; Y = 8'b00010111; // Expected: {'Z': -1794}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110010; Y = 8'b00010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1912,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1794
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000000; Y = 8'b00011101; // Expected: {'Z': -1856}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000000; Y = 8'b00011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1913,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111001; Y = 8'b10011011; // Expected: {'Z': 707}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111001; Y = 8'b10011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1914,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 707
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110010; Y = 8'b10101111; // Expected: {'Z': -4050}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110010; Y = 8'b10101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1915,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011001; Y = 8'b00001110; // Expected: {'Z': 1246}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011001; Y = 8'b00001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1916,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010000; Y = 8'b00111100; // Expected: {'Z': -6720}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010000; Y = 8'b00111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1917,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b01101010; // Expected: {'Z': 1378}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b01101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1918,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1378
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b11111111; // Expected: {'Z': -112}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b11111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1919,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b01101101; // Expected: {'Z': -6431}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b01101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1920,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6431
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010110; Y = 8'b01110100; // Expected: {'Z': -12296}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010110; Y = 8'b01110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1921,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110011; Y = 8'b11000110; // Expected: {'Z': -2958}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110011; Y = 8'b11000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1922,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2958
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011101; Y = 8'b11010000; // Expected: {'Z': 4752}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011101; Y = 8'b11010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1923,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4752
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b10111010; // Expected: {'Z': 4760}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b10111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1924,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101000; Y = 8'b11110011; // Expected: {'Z': -520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101000; Y = 8'b11110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1925,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110010; Y = 8'b11100110; // Expected: {'Z': -2964}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110010; Y = 8'b11100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1926,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2964
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011111; Y = 8'b00010110; // Expected: {'Z': 682}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011111; Y = 8'b00010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1927,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 682
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011100; Y = 8'b11101011; // Expected: {'Z': 756}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011100; Y = 8'b11101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1928,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110000; Y = 8'b11101101; // Expected: {'Z': 1520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110000; Y = 8'b11101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1929,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111110; Y = 8'b00101110; // Expected: {'Z': 2852}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111110; Y = 8'b00101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1930,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2852
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b11001010; // Expected: {'Z': -3996}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b11001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1931,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3996
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000101; Y = 8'b11100110; // Expected: {'Z': -130}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000101; Y = 8'b11100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1932,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110000; Y = 8'b10101001; // Expected: {'Z': -4176}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110000; Y = 8'b10101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1933,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111010; Y = 8'b01001000; // Expected: {'Z': 4176}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111010; Y = 8'b01001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1934,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000001; Y = 8'b01010010; // Expected: {'Z': -5166}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000001; Y = 8'b01010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1935,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011011; Y = 8'b11011011; // Expected: {'Z': -999}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011011; Y = 8'b11011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1936,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -999
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011011; Y = 8'b00010100; // Expected: {'Z': -740}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011011; Y = 8'b00010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1937,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -740
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011010; Y = 8'b11011001; // Expected: {'Z': 3978}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011010; Y = 8'b11011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1938,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3978
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000001; Y = 8'b11101011; // Expected: {'Z': -21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000001; Y = 8'b11101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1939,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001011; Y = 8'b00001001; // Expected: {'Z': -477}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001011; Y = 8'b00001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1940,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -477
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000100; Y = 8'b01110011; // Expected: {'Z': -14260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000100; Y = 8'b01110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1941,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -14260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000111; Y = 8'b11011100; // Expected: {'Z': -252}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000111; Y = 8'b11011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1942,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b11011010; // Expected: {'Z': -342}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b11011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1943,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -342
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011001; Y = 8'b11101011; // Expected: {'Z': -525}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011001; Y = 8'b11101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1944,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -525
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111000; Y = 8'b10000010; // Expected: {'Z': 9072}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111000; Y = 8'b10000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1945,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9072
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100111; Y = 8'b10001000; // Expected: {'Z': 10680}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100111; Y = 8'b10001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1946,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001011; Y = 8'b11010011; // Expected: {'Z': 5265}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001011; Y = 8'b11010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1947,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5265
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111100; Y = 8'b01010001; // Expected: {'Z': 4860}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111100; Y = 8'b01010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1948,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4860
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101011; Y = 8'b10001100; // Expected: {'Z': -4988}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101011; Y = 8'b10001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1949,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4988
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011110; Y = 8'b01011010; // Expected: {'Z': -8820}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011110; Y = 8'b01011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1950,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100010; Y = 8'b01010000; // Expected: {'Z': 7840}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100010; Y = 8'b01010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1951,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000100; Y = 8'b01001010; // Expected: {'Z': -9176}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000100; Y = 8'b01001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1952,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b01011100; // Expected: {'Z': 11316}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b01011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1953,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11316
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010111; Y = 8'b00111000; // Expected: {'Z': 4872}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010111; Y = 8'b00111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1954,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4872
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001100; Y = 8'b01101111; // Expected: {'Z': -12876}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001100; Y = 8'b01101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1955,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12876
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110000; Y = 8'b00000110; // Expected: {'Z': -96}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110000; Y = 8'b00000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1956,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011110; Y = 8'b01010111; // Expected: {'Z': 2610}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011110; Y = 8'b01010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1957,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2610
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011001; Y = 8'b10100010; // Expected: {'Z': -8366}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011001; Y = 8'b10100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1958,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8366
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111001; Y = 8'b11100001; // Expected: {'Z': 217}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111001; Y = 8'b11100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1959,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111101; Y = 8'b00101111; // Expected: {'Z': -141}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111101; Y = 8'b00101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1960,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100111; Y = 8'b00000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100111; Y = 8'b00000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1961,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b01000010; // Expected: {'Z': -3696}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b01000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1962,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3696
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101111; Y = 8'b10001111; // Expected: {'Z': -12543}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101111; Y = 8'b10001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1963,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12543
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100110; Y = 8'b10100011; // Expected: {'Z': -3534}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100110; Y = 8'b10100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1964,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3534
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101110; Y = 8'b10101001; // Expected: {'Z': -4002}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101110; Y = 8'b10101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1965,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4002
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010101; Y = 8'b00001100; // Expected: {'Z': -516}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010101; Y = 8'b00001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1966,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -516
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100011; Y = 8'b01000011; // Expected: {'Z': -1943}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100011; Y = 8'b01000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1967,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1943
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111111; Y = 8'b10111000; // Expected: {'Z': -9144}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111111; Y = 8'b10111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1968,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b00100010; // Expected: {'Z': 3502}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b00100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1969,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3502
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111011; Y = 8'b11110110; // Expected: {'Z': 50}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111011; Y = 8'b11110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1970,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000111; Y = 8'b00000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000111; Y = 8'b00000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1971,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000000; Y = 8'b00101111; // Expected: {'Z': -6016}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000000; Y = 8'b00101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1972,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b01001100; // Expected: {'Z': -5168}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b01001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1973,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b10111010; // Expected: {'Z': -2520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b10111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1974,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101000; Y = 8'b01101101; // Expected: {'Z': -2616}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101000; Y = 8'b01101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1975,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2616
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101000; Y = 8'b11111000; // Expected: {'Z': 192}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101000; Y = 8'b11111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1976,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101001; Y = 8'b10111001; // Expected: {'Z': 1633}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101001; Y = 8'b10111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1977,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1633
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100011; Y = 8'b10101001; // Expected: {'Z': 8091}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100011; Y = 8'b10101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1978,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8091
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001011; Y = 8'b01001010; // Expected: {'Z': 814}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001011; Y = 8'b01001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1979,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 814
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110101; Y = 8'b11001101; // Expected: {'Z': 3825}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110101; Y = 8'b11001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1980,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3825
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010011; Y = 8'b10101010; // Expected: {'Z': 3870}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010011; Y = 8'b10101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1981,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3870
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001100; Y = 8'b01111011; // Expected: {'Z': -6396}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001100; Y = 8'b01111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1982,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6396
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100111; Y = 8'b01000010; // Expected: {'Z': -5874}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100111; Y = 8'b01000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1983,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5874
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110011; Y = 8'b10111011; // Expected: {'Z': -7935}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110011; Y = 8'b10111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1984,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7935
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111110; Y = 8'b11101000; // Expected: {'Z': 1584}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111110; Y = 8'b11101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1985,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1584
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110100; Y = 8'b01110011; // Expected: {'Z': -8740}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110100; Y = 8'b01110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1986,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8740
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111100; Y = 8'b00111111; // Expected: {'Z': 3780}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111100; Y = 8'b00111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1987,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111011; Y = 8'b00100010; // Expected: {'Z': -170}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111011; Y = 8'b00100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1988,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110011; Y = 8'b10010010; // Expected: {'Z': 8470}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110011; Y = 8'b10010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1989,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8470
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110111; Y = 8'b00101110; // Expected: {'Z': 2530}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110111; Y = 8'b00101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1990,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2530
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100100; Y = 8'b11001100; // Expected: {'Z': 4784}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100100; Y = 8'b11001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1991,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111001; Y = 8'b10110000; // Expected: {'Z': 560}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111001; Y = 8'b10110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1992,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111100; Y = 8'b11001111; // Expected: {'Z': -2940}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111100; Y = 8'b11001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1993,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2940
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100110; Y = 8'b11000110; // Expected: {'Z': 5220}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100110; Y = 8'b11000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1994,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111101; Y = 8'b10011011; // Expected: {'Z': 303}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111101; Y = 8'b10011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1995,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 303
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110000; Y = 8'b11111001; // Expected: {'Z': 560}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110000; Y = 8'b11111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1996,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111110; Y = 8'b10101100; // Expected: {'Z': -5208}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111110; Y = 8'b10101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1997,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111111; Y = 8'b00111001; // Expected: {'Z': -57}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111111; Y = 8'b00111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1998,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110101; Y = 8'b10011111; // Expected: {'Z': -5141}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110101; Y = 8'b10011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 1999,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010011; Y = 8'b01000010; // Expected: {'Z': -7194}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010011; Y = 8'b01000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2000,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7194
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100000; Y = 8'b00001001; // Expected: {'Z': -864}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100000; Y = 8'b00001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2001,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -864
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111111; Y = 8'b01000000; // Expected: {'Z': -4160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111111; Y = 8'b01000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2002,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b00000001; // Expected: {'Z': 74}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b00000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2003,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101011; Y = 8'b11001001; // Expected: {'Z': 1155}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101011; Y = 8'b11001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2004,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010001; Y = 8'b01100100; // Expected: {'Z': 1700}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010001; Y = 8'b01100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2005,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011100; Y = 8'b01110101; // Expected: {'Z': 3276}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011100; Y = 8'b01110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2006,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3276
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110001; Y = 8'b11001001; // Expected: {'Z': -2695}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110001; Y = 8'b11001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2007,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2695
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111000; Y = 8'b00001011; // Expected: {'Z': 1320}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111000; Y = 8'b00001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2008,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110011; Y = 8'b01100001; // Expected: {'Z': 4947}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110011; Y = 8'b01100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2009,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4947
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011001; Y = 8'b01010000; // Expected: {'Z': -8240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011001; Y = 8'b01010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2010,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111111; Y = 8'b11011101; // Expected: {'Z': -4445}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111111; Y = 8'b11011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2011,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4445
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011100; Y = 8'b10011111; // Expected: {'Z': 9700}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011100; Y = 8'b10011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2012,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001011; Y = 8'b11111111; // Expected: {'Z': 117}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001011; Y = 8'b11111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2013,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b10100011; // Expected: {'Z': 2604}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b10100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2014,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2604
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100010; Y = 8'b11110101; // Expected: {'Z': 330}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100010; Y = 8'b11110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2015,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 330
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011100; Y = 8'b10111001; // Expected: {'Z': 7100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011100; Y = 8'b10111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2016,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001100; Y = 8'b01011000; // Expected: {'Z': -4576}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001100; Y = 8'b01011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2017,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111001; Y = 8'b00110001; // Expected: {'Z': -3479}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111001; Y = 8'b00110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2018,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3479
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b10100110; // Expected: {'Z': 2520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b10100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2019,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b11110011; // Expected: {'Z': -702}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b11110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2020,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -702
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100011; Y = 8'b01101010; // Expected: {'Z': 10494}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100011; Y = 8'b01101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2021,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10494
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011000; Y = 8'b11101010; // Expected: {'Z': 880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011000; Y = 8'b11101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2022,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000011; Y = 8'b11000100; // Expected: {'Z': 7500}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000011; Y = 8'b11000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2023,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101110; Y = 8'b10011101; // Expected: {'Z': -10890}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101110; Y = 8'b10011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2024,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10890
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b00010101; // Expected: {'Z': 2016}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b00010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2025,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011010; Y = 8'b11101001; // Expected: {'Z': -598}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011010; Y = 8'b11101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2026,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -598
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010101; Y = 8'b00110010; // Expected: {'Z': 4250}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010101; Y = 8'b00110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2027,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101111; Y = 8'b01001000; // Expected: {'Z': -1224}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101111; Y = 8'b01001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2028,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b10000101; // Expected: {'Z': -3567}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b10000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2029,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3567
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000000; Y = 8'b11011010; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000000; Y = 8'b11011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2030,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b00110111; // Expected: {'Z': -3245}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b00110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2031,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001100; Y = 8'b01011000; // Expected: {'Z': -10208}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001100; Y = 8'b01011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2032,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001010; Y = 8'b10011110; // Expected: {'Z': -980}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001010; Y = 8'b10011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2033,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011010; Y = 8'b00111100; // Expected: {'Z': 5400}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011010; Y = 8'b00111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2034,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011000; Y = 8'b10011011; // Expected: {'Z': 10504}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011000; Y = 8'b10011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2035,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101010; Y = 8'b01000010; // Expected: {'Z': -1452}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101010; Y = 8'b01000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2036,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1452
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b10000000; // Expected: {'Z': 7168}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b10000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2037,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001111; Y = 8'b00100111; // Expected: {'Z': -1911}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001111; Y = 8'b00100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2038,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1911
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000100; Y = 8'b01010011; // Expected: {'Z': -4980}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000100; Y = 8'b01010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2039,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110010; Y = 8'b11100100; // Expected: {'Z': 392}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110010; Y = 8'b11100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2040,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110011; Y = 8'b10010011; // Expected: {'Z': -12535}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110011; Y = 8'b10010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2041,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12535
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111011; Y = 8'b10011001; // Expected: {'Z': 7107}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111011; Y = 8'b10011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2042,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110100; Y = 8'b01101001; // Expected: {'Z': -1260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110100; Y = 8'b01101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2043,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b00101100; // Expected: {'Z': -2992}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b00101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2044,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2992
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101000; Y = 8'b01111111; // Expected: {'Z': 13208}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101000; Y = 8'b01111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2045,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 13208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b11101011; // Expected: {'Z': -462}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b11101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2046,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111000; Y = 8'b00011100; // Expected: {'Z': -2016}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111000; Y = 8'b00011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2047,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b00101000; // Expected: {'Z': -2040}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b00101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2048,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000101; Y = 8'b01011100; // Expected: {'Z': 6348}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000101; Y = 8'b01011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2049,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6348
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010000; Y = 8'b10101100; // Expected: {'Z': -6720}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010000; Y = 8'b10101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2050,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110101; Y = 8'b01110011; // Expected: {'Z': 13455}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110101; Y = 8'b01110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2051,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 13455
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010110; Y = 8'b11011110; // Expected: {'Z': 3604}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010110; Y = 8'b11011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2052,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3604
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011111; Y = 8'b11111101; // Expected: {'Z': 99}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011111; Y = 8'b11111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2053,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b01111110; // Expected: {'Z': 2394}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b01111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2054,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2394
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010010; Y = 8'b10100010; // Expected: {'Z': -1692}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010010; Y = 8'b10100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2055,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1692
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b10011111; // Expected: {'Z': -1261}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b10011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2056,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1261
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111100; Y = 8'b00011111; // Expected: {'Z': 1860}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111100; Y = 8'b00011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2057,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1860
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001100; Y = 8'b10011110; // Expected: {'Z': 5096}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001100; Y = 8'b10011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2058,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5096
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111000; Y = 8'b11001010; // Expected: {'Z': 432}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111000; Y = 8'b11001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2059,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100011; Y = 8'b11110000; // Expected: {'Z': 464}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100011; Y = 8'b11110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2060,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111110; Y = 8'b10000100; // Expected: {'Z': -15624}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111110; Y = 8'b10000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2061,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -15624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100010; Y = 8'b11001101; // Expected: {'Z': -4998}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100010; Y = 8'b11001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2062,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4998
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111010; Y = 8'b11011000; // Expected: {'Z': 2800}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111010; Y = 8'b11011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2063,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011010; Y = 8'b00101110; // Expected: {'Z': 1196}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011010; Y = 8'b00101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2064,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011000; Y = 8'b01000111; // Expected: {'Z': -7384}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011000; Y = 8'b01000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2065,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7384
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000001; Y = 8'b01011110; // Expected: {'Z': -5922}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000001; Y = 8'b01011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2066,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5922
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101111; Y = 8'b00110001; // Expected: {'Z': 5439}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101111; Y = 8'b00110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2067,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5439
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001100; Y = 8'b11110011; // Expected: {'Z': -156}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001100; Y = 8'b11110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2068,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011011; Y = 8'b01100011; // Expected: {'Z': 9009}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011011; Y = 8'b01100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2069,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9009
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101010; Y = 8'b10101111; // Expected: {'Z': 1782}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101010; Y = 8'b10101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2070,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1782
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111001; Y = 8'b01001001; // Expected: {'Z': 8833}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111001; Y = 8'b01001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2071,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8833
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100100; Y = 8'b01010101; // Expected: {'Z': -7820}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100100; Y = 8'b01010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2072,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111011; Y = 8'b11100111; // Expected: {'Z': 1725}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111011; Y = 8'b11100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2073,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1725
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111000; Y = 8'b00011110; // Expected: {'Z': 1680}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111000; Y = 8'b00011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2074,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b00001011; // Expected: {'Z': 484}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b00001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2075,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 484
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010000; Y = 8'b01011010; // Expected: {'Z': -4320}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010000; Y = 8'b01011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2076,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000100; Y = 8'b10001110; // Expected: {'Z': 6840}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000100; Y = 8'b10001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2077,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011110; Y = 8'b10111100; // Expected: {'Z': 6664}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011110; Y = 8'b10111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2078,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6664
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010111; Y = 8'b11000110; // Expected: {'Z': -5046}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010111; Y = 8'b11000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2079,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5046
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010101; Y = 8'b11111100; // Expected: {'Z': -340}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010101; Y = 8'b11111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2080,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010000; Y = 8'b11001011; // Expected: {'Z': 5936}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010000; Y = 8'b11001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2081,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5936
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110111; Y = 8'b10100000; // Expected: {'Z': -11424}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110111; Y = 8'b10100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2082,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11424
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010101; Y = 8'b01101110; // Expected: {'Z': -11770}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010101; Y = 8'b01101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2083,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11770
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b10100101; // Expected: {'Z': -819}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b10100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2084,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -819
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011110; Y = 8'b10110001; // Expected: {'Z': -7426}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011110; Y = 8'b10110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2085,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7426
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001011; Y = 8'b00111010; // Expected: {'Z': 4350}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001011; Y = 8'b00111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2086,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010000; Y = 8'b11100101; // Expected: {'Z': -2160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010000; Y = 8'b11100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2087,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000011; Y = 8'b10110001; // Expected: {'Z': -5293}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000011; Y = 8'b10110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2088,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5293
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b11001010; // Expected: {'Z': -1134}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b11001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2089,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101100; Y = 8'b00101000; // Expected: {'Z': -800}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101100; Y = 8'b00101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2090,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001011; Y = 8'b00110000; // Expected: {'Z': -2544}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001011; Y = 8'b00110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2091,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2544
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100100; Y = 8'b10000011; // Expected: {'Z': 11500}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100100; Y = 8'b10000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2092,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010101; Y = 8'b00000010; // Expected: {'Z': -86}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010101; Y = 8'b00000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2093,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b01110100; // Expected: {'Z': 4176}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b01110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2094,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b10000101; // Expected: {'Z': -1599}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b10000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2095,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1599
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010001; Y = 8'b10101000; // Expected: {'Z': -7128}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010001; Y = 8'b10101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2096,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110110; Y = 8'b01101001; // Expected: {'Z': 12390}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110110; Y = 8'b01101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2097,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 12390
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010100; Y = 8'b01011001; // Expected: {'Z': 7476}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010100; Y = 8'b01011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2098,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7476
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011011; Y = 8'b11111110; // Expected: {'Z': 202}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011011; Y = 8'b11111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2099,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011110; Y = 8'b10000011; // Expected: {'Z': -3750}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011110; Y = 8'b10000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2100,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100001; Y = 8'b01011111; // Expected: {'Z': 3135}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100001; Y = 8'b01011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2101,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010110; Y = 8'b11110010; // Expected: {'Z': -1204}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010110; Y = 8'b11110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2102,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b11001100; // Expected: {'Z': -5824}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b11001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2103,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5824
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001100; Y = 8'b01111101; // Expected: {'Z': -6500}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001100; Y = 8'b01111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2104,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b11010011; // Expected: {'Z': -3960}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b11010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2105,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011100; Y = 8'b00001011; // Expected: {'Z': -396}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011100; Y = 8'b00001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2106,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -396
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011110; Y = 8'b00010000; // Expected: {'Z': 1504}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011110; Y = 8'b00010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2107,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101100; Y = 8'b00011101; // Expected: {'Z': -580}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101100; Y = 8'b00011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2108,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010000; Y = 8'b10010101; // Expected: {'Z': 11984}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010000; Y = 8'b10010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2109,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11984
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b01110001; // Expected: {'Z': 2373}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b01110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2110,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2373
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110011; Y = 8'b00111101; // Expected: {'Z': -793}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110011; Y = 8'b00111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2111,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -793
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010010; Y = 8'b01101001; // Expected: {'Z': -11550}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010010; Y = 8'b01101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2112,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b10111101; // Expected: {'Z': -134}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b10111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2113,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110101; Y = 8'b01000001; // Expected: {'Z': 3445}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110101; Y = 8'b01000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2114,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3445
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b00011000; // Expected: {'Z': 696}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b00011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2115,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 696
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101010; Y = 8'b11110000; // Expected: {'Z': 1376}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101010; Y = 8'b11110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2116,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1376
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101000; Y = 8'b10011000; // Expected: {'Z': -10816}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101000; Y = 8'b10011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2117,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b10001100; // Expected: {'Z': -4176}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b10001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2118,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010111; Y = 8'b10101011; // Expected: {'Z': 8925}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010111; Y = 8'b10101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2119,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8925
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111110; Y = 8'b01011100; // Expected: {'Z': -6072}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111110; Y = 8'b01011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2120,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6072
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b01000000; // Expected: {'Z': 960}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b01000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2121,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111011; Y = 8'b01011001; // Expected: {'Z': -445}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111011; Y = 8'b01011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2122,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -445
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010001; Y = 8'b11111000; // Expected: {'Z': -136}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010001; Y = 8'b11111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2123,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001000; Y = 8'b11000000; // Expected: {'Z': -512}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001000; Y = 8'b11000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2124,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -512
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b10101000; // Expected: {'Z': 5984}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b10101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2125,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5984
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110000; Y = 8'b01100100; // Expected: {'Z': -1600}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110000; Y = 8'b01100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2126,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110011; Y = 8'b01111101; // Expected: {'Z': 14375}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110011; Y = 8'b01111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2127,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 14375
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101001; Y = 8'b01000001; // Expected: {'Z': 2665}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101001; Y = 8'b01000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2128,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2665
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101101; Y = 8'b11101111; // Expected: {'Z': -765}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101101; Y = 8'b11101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2129,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -765
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010001; Y = 8'b10100101; // Expected: {'Z': -7371}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010001; Y = 8'b10100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2130,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7371
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000000; Y = 8'b11111010; // Expected: {'Z': 384}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000000; Y = 8'b11111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2131,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 384
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011011; Y = 8'b10010100; // Expected: {'Z': -2916}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011011; Y = 8'b10010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2132,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2916
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100001; Y = 8'b00011000; // Expected: {'Z': 2328}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100001; Y = 8'b00011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2133,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2328
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110110; Y = 8'b00100111; // Expected: {'Z': -390}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110110; Y = 8'b00100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2134,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -390
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110101; Y = 8'b10001011; // Expected: {'Z': 8775}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110101; Y = 8'b10001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2135,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8775
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100011; Y = 8'b11101000; // Expected: {'Z': 696}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100011; Y = 8'b11101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2136,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 696
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011111; Y = 8'b10100001; // Expected: {'Z': 9215}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011111; Y = 8'b10100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2137,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9215
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b11001000; // Expected: {'Z': 3136}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b11001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2138,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100011; Y = 8'b11101100; // Expected: {'Z': -700}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100011; Y = 8'b11101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2139,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111100; Y = 8'b10111010; // Expected: {'Z': -8680}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111100; Y = 8'b10111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2140,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101101; Y = 8'b10011110; // Expected: {'Z': -10682}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101101; Y = 8'b10011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2141,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10682
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000001; Y = 8'b10100100; // Expected: {'Z': -92}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000001; Y = 8'b10100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2142,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100101; Y = 8'b10001100; // Expected: {'Z': -11716}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100101; Y = 8'b10001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2143,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11716
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101000; Y = 8'b11010100; // Expected: {'Z': -1760}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101000; Y = 8'b11010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2144,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101010; Y = 8'b01001010; // Expected: {'Z': -6364}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101010; Y = 8'b01001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2145,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110101; Y = 8'b01001100; // Expected: {'Z': -5700}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110101; Y = 8'b01001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2146,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100010; Y = 8'b11000110; // Expected: {'Z': -5684}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100010; Y = 8'b11000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2147,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5684
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111110; Y = 8'b01000011; // Expected: {'Z': -134}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111110; Y = 8'b01000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2148,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b10000011; // Expected: {'Z': 8500}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b10000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2149,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001111; Y = 8'b11101100; // Expected: {'Z': -1580}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001111; Y = 8'b11101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2150,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011010; Y = 8'b10011110; // Expected: {'Z': 3724}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011010; Y = 8'b10011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2151,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3724
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111000; Y = 8'b11110010; // Expected: {'Z': -1680}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111000; Y = 8'b11110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2152,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b11000101; // Expected: {'Z': -885}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b11000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2153,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -885
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110100; Y = 8'b11011101; // Expected: {'Z': -4060}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110100; Y = 8'b11011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2154,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100110; Y = 8'b11111101; // Expected: {'Z': -306}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100110; Y = 8'b11111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2155,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -306
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101111; Y = 8'b00000001; // Expected: {'Z': -81}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101111; Y = 8'b00000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2156,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000001; Y = 8'b01001010; // Expected: {'Z': -4662}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000001; Y = 8'b01001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2157,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4662
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101101; Y = 8'b00101000; // Expected: {'Z': -3320}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101101; Y = 8'b00101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2158,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000000; Y = 8'b10000010; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000000; Y = 8'b10000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2159,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010001; Y = 8'b10100101; // Expected: {'Z': 4277}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010001; Y = 8'b10100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2160,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4277
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100010; Y = 8'b11001001; // Expected: {'Z': 1650}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100010; Y = 8'b11001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2161,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011010; Y = 8'b01010101; // Expected: {'Z': 2210}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011010; Y = 8'b01010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2162,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010011; Y = 8'b00100111; // Expected: {'Z': -4251}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010011; Y = 8'b00100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2163,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001111; Y = 8'b11100110; // Expected: {'Z': -2054}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001111; Y = 8'b11100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2164,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2054
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000010; Y = 8'b00100101; // Expected: {'Z': 2442}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000010; Y = 8'b00100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2165,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2442
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010011; Y = 8'b00001100; // Expected: {'Z': 996}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010011; Y = 8'b00001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2166,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 996
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101101; Y = 8'b00101100; // Expected: {'Z': 1980}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101101; Y = 8'b00101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2167,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111001; Y = 8'b11101011; // Expected: {'Z': -2541}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111001; Y = 8'b11101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2168,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2541
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011010; Y = 8'b10001001; // Expected: {'Z': -10710}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011010; Y = 8'b10001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2169,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10710
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b10000110; // Expected: {'Z': 7198}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b10000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2170,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b10011011; // Expected: {'Z': 5959}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b10011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2171,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5959
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000001; Y = 8'b10000111; // Expected: {'Z': 15367}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000001; Y = 8'b10000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2172,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 15367
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b01110111; // Expected: {'Z': 12257}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b01110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2173,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 12257
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b00000110; // Expected: {'Z': -504}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b00000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2174,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b10001011; // Expected: {'Z': -234}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b10001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2175,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101011; Y = 8'b01010111; // Expected: {'Z': 3741}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101011; Y = 8'b01010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2176,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3741
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010101; Y = 8'b00100101; // Expected: {'Z': 3145}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010101; Y = 8'b00100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2177,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001111; Y = 8'b10010110; // Expected: {'Z': -8374}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001111; Y = 8'b10010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2178,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8374
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b00111100; // Expected: {'Z': 6180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b00111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2179,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100000; Y = 8'b11101101; // Expected: {'Z': 608}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100000; Y = 8'b11101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2180,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 608
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000000; Y = 8'b00000001; // Expected: {'Z': -128}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000000; Y = 8'b00000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2181,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b00110000; // Expected: {'Z': 3552}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b00110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2182,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110110; Y = 8'b00010000; // Expected: {'Z': 1888}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110110; Y = 8'b00010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2183,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100110; Y = 8'b01101101; // Expected: {'Z': 11118}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100110; Y = 8'b01101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2184,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000110; Y = 8'b00000100; // Expected: {'Z': -488}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000110; Y = 8'b00000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2185,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110000; Y = 8'b10100011; // Expected: {'Z': 1488}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110000; Y = 8'b10100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2186,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111101; Y = 8'b01100101; // Expected: {'Z': -6767}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111101; Y = 8'b01100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2187,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6767
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000001; Y = 8'b00111010; // Expected: {'Z': 58}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000001; Y = 8'b00111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2188,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011100; Y = 8'b11111011; // Expected: {'Z': -140}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011100; Y = 8'b11111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2189,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101001; Y = 8'b01000101; // Expected: {'Z': 7245}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101001; Y = 8'b01000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2190,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000000; Y = 8'b10010000; // Expected: {'Z': 14336}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000000; Y = 8'b10010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2191,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 14336
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011100; Y = 8'b10111010; // Expected: {'Z': 7000}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011100; Y = 8'b10111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2192,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110010; Y = 8'b00100010; // Expected: {'Z': -2652}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110010; Y = 8'b00100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2193,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2652
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100110; Y = 8'b11100000; // Expected: {'Z': -1216}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100110; Y = 8'b11100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2194,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000110; Y = 8'b01110000; // Expected: {'Z': -13664}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000110; Y = 8'b01110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2195,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -13664
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011010; Y = 8'b01100011; // Expected: {'Z': -3762}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011010; Y = 8'b01100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2196,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3762
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101110; Y = 8'b00100100; // Expected: {'Z': -648}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101110; Y = 8'b00100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2197,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011100; Y = 8'b10011101; // Expected: {'Z': 3564}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011100; Y = 8'b10011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2198,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3564
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011001; Y = 8'b11001101; // Expected: {'Z': 1989}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011001; Y = 8'b11001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2199,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1989
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101011; Y = 8'b01001001; // Expected: {'Z': -1533}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101011; Y = 8'b01001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2200,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1533
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011011; Y = 8'b01001011; // Expected: {'Z': 2025}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011011; Y = 8'b01001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2201,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2025
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b00111101; // Expected: {'Z': 4514}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b00111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2202,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4514
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010000; Y = 8'b10011110; // Expected: {'Z': 10976}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010000; Y = 8'b10011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2203,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10976
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111101; Y = 8'b11111110; // Expected: {'Z': -250}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111101; Y = 8'b11111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2204,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011110; Y = 8'b11100111; // Expected: {'Z': 2450}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011110; Y = 8'b11100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2205,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011100; Y = 8'b10111010; // Expected: {'Z': -6440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011100; Y = 8'b10111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2206,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100010; Y = 8'b01011110; // Expected: {'Z': 3196}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100010; Y = 8'b01011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2207,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111110; Y = 8'b10010001; // Expected: {'Z': 7326}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111110; Y = 8'b10010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2208,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7326
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001000; Y = 8'b10010110; // Expected: {'Z': -848}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001000; Y = 8'b10010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2209,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110100; Y = 8'b10001001; // Expected: {'Z': -6188}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110100; Y = 8'b10001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2210,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111101; Y = 8'b01001011; // Expected: {'Z': -5025}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111101; Y = 8'b01001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2211,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5025
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b11000101; // Expected: {'Z': -354}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b11000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2212,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -354
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000001; Y = 8'b10000111; // Expected: {'Z': 7623}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000001; Y = 8'b10000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2213,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7623
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b10000100; // Expected: {'Z': -744}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b10000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2214,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -744
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101101; Y = 8'b01101110; // Expected: {'Z': -2090}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101101; Y = 8'b01101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2215,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2090
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111000; Y = 8'b10011010; // Expected: {'Z': -12240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111000; Y = 8'b10011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2216,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010001; Y = 8'b00111111; // Expected: {'Z': -2961}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010001; Y = 8'b00111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2217,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2961
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110001; Y = 8'b10100010; // Expected: {'Z': -4606}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110001; Y = 8'b10100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2218,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4606
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b11001110; // Expected: {'Z': -4400}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b11001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2219,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101000; Y = 8'b00010001; // Expected: {'Z': 680}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101000; Y = 8'b00010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2220,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b10000001; // Expected: {'Z': -15621}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b10000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2221,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -15621
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b01001101; // Expected: {'Z': 3003}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b01001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2222,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3003
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101000; Y = 8'b10110111; // Expected: {'Z': -2920}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101000; Y = 8'b10110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2223,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010110; Y = 8'b10110101; // Expected: {'Z': 3150}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010110; Y = 8'b10110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2224,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011101; Y = 8'b00000101; // Expected: {'Z': 465}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011101; Y = 8'b00000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2225,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 465
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111111; Y = 8'b10010011; // Expected: {'Z': 109}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111111; Y = 8'b10010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2226,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 109
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110000; Y = 8'b00110010; // Expected: {'Z': -800}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110000; Y = 8'b00110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2227,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101101; Y = 8'b00000100; // Expected: {'Z': 436}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101101; Y = 8'b00000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2228,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 436
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100000; Y = 8'b00001011; // Expected: {'Z': -1056}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100000; Y = 8'b00001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2229,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1056
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010011; Y = 8'b00011101; // Expected: {'Z': -3161}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010011; Y = 8'b00011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2230,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3161
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001011; Y = 8'b00100110; // Expected: {'Z': -2014}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001011; Y = 8'b00100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2231,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2014
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001001; Y = 8'b01011101; // Expected: {'Z': 6789}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001001; Y = 8'b01011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2232,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6789
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b11000011; // Expected: {'Z': 5124}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b11000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2233,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101010; Y = 8'b10101100; // Expected: {'Z': 7224}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101010; Y = 8'b10101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2234,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100001; Y = 8'b10100110; // Expected: {'Z': -2970}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100001; Y = 8'b10100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2235,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2970
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111011; Y = 8'b01111111; // Expected: {'Z': -8763}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111011; Y = 8'b01111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2236,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8763
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101011; Y = 8'b00000010; // Expected: {'Z': -170}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101011; Y = 8'b00000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2237,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000001; Y = 8'b00100110; // Expected: {'Z': -2394}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000001; Y = 8'b00100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2238,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2394
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100110; Y = 8'b10110100; // Expected: {'Z': -2888}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100110; Y = 8'b10110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2239,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100111; Y = 8'b11100010; // Expected: {'Z': 2670}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100111; Y = 8'b11100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2240,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2670
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100100; Y = 8'b11110011; // Expected: {'Z': 1196}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100100; Y = 8'b11110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2241,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101111; Y = 8'b10110101; // Expected: {'Z': -8325}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101111; Y = 8'b10110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2242,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8325
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001100; Y = 8'b01100011; // Expected: {'Z': -5148}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001100; Y = 8'b01100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2243,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001011; Y = 8'b01101011; // Expected: {'Z': -5671}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001011; Y = 8'b01101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2244,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5671
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000011; Y = 8'b11100100; // Expected: {'Z': -84}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000011; Y = 8'b11100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2245,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011010; Y = 8'b01000010; // Expected: {'Z': 5940}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011010; Y = 8'b01000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2246,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5940
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111010; Y = 8'b01000010; // Expected: {'Z': -396}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111010; Y = 8'b01000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2247,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -396
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000000; Y = 8'b01011001; // Expected: {'Z': -11392}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000000; Y = 8'b01011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2248,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110011; Y = 8'b01100001; // Expected: {'Z': -1261}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110011; Y = 8'b01100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2249,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1261
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110001; Y = 8'b01000011; // Expected: {'Z': -1005}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110001; Y = 8'b01000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2250,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1005
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b00011111; // Expected: {'Z': 403}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b00011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2251,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 403
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100000; Y = 8'b00111100; // Expected: {'Z': 1920}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100000; Y = 8'b00111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2252,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b00010101; // Expected: {'Z': 1134}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b00010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2253,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100000; Y = 8'b10110100; // Expected: {'Z': 7296}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100000; Y = 8'b10110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2254,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111111; Y = 8'b10111101; // Expected: {'Z': -4221}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111111; Y = 8'b10111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2255,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b11110001; // Expected: {'Z': 1260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b11110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2256,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000010; Y = 8'b10000111; // Expected: {'Z': -7986}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000010; Y = 8'b10000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2257,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7986
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000010; Y = 8'b10000100; // Expected: {'Z': 7688}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000010; Y = 8'b10000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2258,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7688
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010101; Y = 8'b00000010; // Expected: {'Z': -86}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010101; Y = 8'b00000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2259,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101001; Y = 8'b11100110; // Expected: {'Z': -2730}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101001; Y = 8'b11100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2260,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2730
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000101; Y = 8'b11111011; // Expected: {'Z': 615}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000101; Y = 8'b11111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2261,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 615
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b10000011; // Expected: {'Z': -6750}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b10000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2262,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111010; Y = 8'b00110001; // Expected: {'Z': 2842}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111010; Y = 8'b00110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2263,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2842
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010111; Y = 8'b00011100; // Expected: {'Z': -1148}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010111; Y = 8'b00011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2264,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100101; Y = 8'b11101001; // Expected: {'Z': 621}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100101; Y = 8'b11101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2265,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 621
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010000; Y = 8'b10110010; // Expected: {'Z': -6240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010000; Y = 8'b10110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2266,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110110; Y = 8'b00000010; // Expected: {'Z': 236}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110110; Y = 8'b00000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2267,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010010; Y = 8'b11011101; // Expected: {'Z': 3850}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010010; Y = 8'b11011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2268,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3850
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101101; Y = 8'b00100110; // Expected: {'Z': -722}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101101; Y = 8'b00100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2269,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -722
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110100; Y = 8'b10101110; // Expected: {'Z': -9512}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110100; Y = 8'b10101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2270,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9512
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011110; Y = 8'b00111010; // Expected: {'Z': -1972}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011110; Y = 8'b00111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2271,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1972
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110001; Y = 8'b11101100; // Expected: {'Z': 300}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110001; Y = 8'b11101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2272,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011110; Y = 8'b00010010; // Expected: {'Z': 1692}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011110; Y = 8'b00010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2273,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1692
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101110; Y = 8'b10101111; // Expected: {'Z': -8910}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101110; Y = 8'b10101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2274,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8910
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011000; Y = 8'b00011011; // Expected: {'Z': -1080}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011000; Y = 8'b00011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2275,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111101; Y = 8'b01101011; // Expected: {'Z': -321}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111101; Y = 8'b01101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2276,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -321
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001100; Y = 8'b01001101; // Expected: {'Z': 924}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001100; Y = 8'b01001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2277,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 924
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b10111111; // Expected: {'Z': -4680}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b10111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2278,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000000; Y = 8'b11110011; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000000; Y = 8'b11110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2279,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100000; Y = 8'b10100110; // Expected: {'Z': 2880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100000; Y = 8'b10100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2280,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100000; Y = 8'b10111010; // Expected: {'Z': 2240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100000; Y = 8'b10111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2281,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100110; Y = 8'b00101000; // Expected: {'Z': 1520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100110; Y = 8'b00101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2282,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011010; Y = 8'b11001001; // Expected: {'Z': -1430}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011010; Y = 8'b11001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2283,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000011; Y = 8'b10000101; // Expected: {'Z': -369}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000011; Y = 8'b10000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2284,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -369
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100011; Y = 8'b01110101; // Expected: {'Z': 11583}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100011; Y = 8'b01110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2285,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11583
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010010; Y = 8'b01100110; // Expected: {'Z': 1836}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010010; Y = 8'b01100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2286,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1836
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010010; Y = 8'b10010110; // Expected: {'Z': 11660}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010010; Y = 8'b10010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2287,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000010; Y = 8'b00011101; // Expected: {'Z': -3654}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000010; Y = 8'b00011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2288,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3654
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011100; Y = 8'b01010101; // Expected: {'Z': 7820}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011100; Y = 8'b01010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2289,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101010; Y = 8'b10111101; // Expected: {'Z': 1474}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101010; Y = 8'b10111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2290,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1474
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100001; Y = 8'b11110001; // Expected: {'Z': -1455}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100001; Y = 8'b11110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2291,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1455
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001001; Y = 8'b11110011; // Expected: {'Z': 1547}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001001; Y = 8'b11110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2292,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1547
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011001; Y = 8'b00011100; // Expected: {'Z': 700}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011001; Y = 8'b00011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2293,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011100; Y = 8'b00001011; // Expected: {'Z': -1100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011100; Y = 8'b00001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2294,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101111; Y = 8'b11110011; // Expected: {'Z': -1443}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101111; Y = 8'b11110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2295,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1443
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101000; Y = 8'b11011111; // Expected: {'Z': -3432}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101000; Y = 8'b11011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2296,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010101; Y = 8'b10101110; // Expected: {'Z': 8774}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010101; Y = 8'b10101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2297,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8774
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111111; Y = 8'b10111101; // Expected: {'Z': 4355}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111111; Y = 8'b10111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2298,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4355
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110010; Y = 8'b10010001; // Expected: {'Z': -12654}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110010; Y = 8'b10010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2299,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12654
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110111; Y = 8'b11001011; // Expected: {'Z': 477}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110111; Y = 8'b11001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2300,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 477
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000000; Y = 8'b11111011; // Expected: {'Z': 640}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000000; Y = 8'b11111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2301,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001100; Y = 8'b00001101; // Expected: {'Z': 156}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001100; Y = 8'b00001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2302,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100110; Y = 8'b01011011; // Expected: {'Z': -2366}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100110; Y = 8'b01011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2303,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2366
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111000; Y = 8'b11010110; // Expected: {'Z': -2352}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111000; Y = 8'b11010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2304,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b10000101; // Expected: {'Z': 6273}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b10000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2305,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6273
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000000; Y = 8'b00010001; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000000; Y = 8'b00010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2306,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000011; Y = 8'b00001101; // Expected: {'Z': -1625}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000011; Y = 8'b00001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2307,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1625
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b11110010; // Expected: {'Z': -756}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b11110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2308,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000101; Y = 8'b01100100; // Expected: {'Z': -12300}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000101; Y = 8'b01100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2309,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110111; Y = 8'b10011010; // Expected: {'Z': 918}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110111; Y = 8'b10011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2310,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 918
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011100; Y = 8'b01111101; // Expected: {'Z': 11500}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011100; Y = 8'b01111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2311,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b00100010; // Expected: {'Z': 204}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b00100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2312,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000101; Y = 8'b11100011; // Expected: {'Z': -2001}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000101; Y = 8'b11100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2313,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2001
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b10011001; // Expected: {'Z': -3708}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b10011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2314,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3708
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001011; Y = 8'b11000110; // Expected: {'Z': -638}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001011; Y = 8'b11000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2315,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -638
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010011; Y = 8'b11000110; // Expected: {'Z': 6322}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010011; Y = 8'b11000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2316,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6322
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111101; Y = 8'b01001010; // Expected: {'Z': -4958}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111101; Y = 8'b01001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2317,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4958
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011011; Y = 8'b01001100; // Expected: {'Z': 2052}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011011; Y = 8'b01001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2318,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2052
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b10100110; // Expected: {'Z': -11070}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b10100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2319,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11070
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101010; Y = 8'b10011101; // Expected: {'Z': -4158}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101010; Y = 8'b10011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2320,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4158
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110001; Y = 8'b10011000; // Expected: {'Z': -5096}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110001; Y = 8'b10011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2321,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5096
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101110; Y = 8'b10110100; // Expected: {'Z': -3496}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101110; Y = 8'b10110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2322,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b11110001; // Expected: {'Z': 1260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b11110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2323,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011011; Y = 8'b10110111; // Expected: {'Z': -1971}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011011; Y = 8'b10110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2324,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1971
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110110; Y = 8'b00001000; // Expected: {'Z': -592}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110110; Y = 8'b00001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2325,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -592
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100010; Y = 8'b01011100; // Expected: {'Z': -8648}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100010; Y = 8'b01011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2326,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011111; Y = 8'b11111010; // Expected: {'Z': 582}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011111; Y = 8'b11111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2327,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 582
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110010; Y = 8'b01011001; // Expected: {'Z': 10146}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110010; Y = 8'b01011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2328,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110111; Y = 8'b11010000; // Expected: {'Z': -2640}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110111; Y = 8'b11010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2329,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b00000011; // Expected: {'Z': 264}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b00000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2330,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000100; Y = 8'b00100010; // Expected: {'Z': 136}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000100; Y = 8'b00100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2331,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b01100110; // Expected: {'Z': -5712}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b01100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2332,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5712
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110110; Y = 8'b00001001; // Expected: {'Z': -90}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110110; Y = 8'b00001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2333,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110011; Y = 8'b10001011; // Expected: {'Z': 1521}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110011; Y = 8'b10001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2334,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1521
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000011; Y = 8'b00111000; // Expected: {'Z': 168}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000011; Y = 8'b00111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2335,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001100; Y = 8'b10111010; // Expected: {'Z': -5320}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001100; Y = 8'b10111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2336,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b00000011; // Expected: {'Z': 132}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b00000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2337,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b00100010; // Expected: {'Z': 1598}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b00100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2338,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1598
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101000; Y = 8'b10011000; // Expected: {'Z': -10816}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101000; Y = 8'b10011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2339,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110111; Y = 8'b11000111; // Expected: {'Z': -6783}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110111; Y = 8'b11000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2340,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6783
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011001; Y = 8'b11110101; // Expected: {'Z': -275}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011001; Y = 8'b11110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2341,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -275
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100111; Y = 8'b10010000; // Expected: {'Z': 9968}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100111; Y = 8'b10010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2342,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9968
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011011; Y = 8'b10000011; // Expected: {'Z': -3375}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011011; Y = 8'b10000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2343,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3375
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110111; Y = 8'b10101010; // Expected: {'Z': 6278}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110111; Y = 8'b10101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2344,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6278
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111110; Y = 8'b01111010; // Expected: {'Z': 15372}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111110; Y = 8'b01111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2345,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 15372
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b01100110; // Expected: {'Z': -6936}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b01100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2346,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6936
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011111; Y = 8'b01010011; // Expected: {'Z': -2739}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011111; Y = 8'b01010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2347,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2739
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b11010101; // Expected: {'Z': -258}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b11010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2348,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -258
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000000; Y = 8'b01001101; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000000; Y = 8'b01001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2349,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010001; Y = 8'b01000011; // Expected: {'Z': 1139}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010001; Y = 8'b01000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2350,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1139
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010010; Y = 8'b01100111; // Expected: {'Z': -11330}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010010; Y = 8'b01100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2351,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11330
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111010; Y = 8'b10111100; // Expected: {'Z': -3944}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111010; Y = 8'b10111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2352,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b00101011; // Expected: {'Z': -4773}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b00101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2353,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4773
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b01101110; // Expected: {'Z': 660}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b01101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2354,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110000; Y = 8'b10000101; // Expected: {'Z': 9840}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110000; Y = 8'b10000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2355,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001100; Y = 8'b11011101; // Expected: {'Z': 1820}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001100; Y = 8'b11011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2356,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011101; Y = 8'b01011000; // Expected: {'Z': -8712}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011101; Y = 8'b01011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2357,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8712
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011110; Y = 8'b10100000; // Expected: {'Z': 9408}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011110; Y = 8'b10100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2358,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b01010111; // Expected: {'Z': 1827}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b01010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2359,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1827
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010011; Y = 8'b00000110; // Expected: {'Z': -654}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010011; Y = 8'b00000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2360,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -654
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010001; Y = 8'b10010010; // Expected: {'Z': 5170}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010001; Y = 8'b10010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2361,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000111; Y = 8'b11100110; // Expected: {'Z': -1846}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000111; Y = 8'b11100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2362,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1846
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110001; Y = 8'b10100000; // Expected: {'Z': -10848}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110001; Y = 8'b10100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2363,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000000; Y = 8'b01110101; // Expected: {'Z': -14976}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000000; Y = 8'b01110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2364,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -14976
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b01001010; // Expected: {'Z': 7622}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b01001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2365,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7622
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101011; Y = 8'b00010110; // Expected: {'Z': -462}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101011; Y = 8'b00010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2366,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111000; Y = 8'b11101001; // Expected: {'Z': 1656}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111000; Y = 8'b11101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2367,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1656
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010110; Y = 8'b01110000; // Expected: {'Z': 9632}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010110; Y = 8'b01110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2368,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9632
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111010; Y = 8'b00011010; // Expected: {'Z': 1508}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111010; Y = 8'b00011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2369,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1508
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110000; Y = 8'b01111101; // Expected: {'Z': -2000}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110000; Y = 8'b01111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2370,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010110; Y = 8'b11011001; // Expected: {'Z': -3354}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010110; Y = 8'b11011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2371,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3354
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100010; Y = 8'b00101111; // Expected: {'Z': 1598}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100010; Y = 8'b00101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2372,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1598
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b01011011; // Expected: {'Z': 182}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b01011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2373,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011001; Y = 8'b00100101; // Expected: {'Z': -3811}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011001; Y = 8'b00100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2374,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3811
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101010; Y = 8'b11110010; // Expected: {'Z': -588}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101010; Y = 8'b11110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2375,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -588
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111111; Y = 8'b10110110; // Expected: {'Z': -9398}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111111; Y = 8'b10110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2376,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9398
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000011; Y = 8'b00011010; // Expected: {'Z': 1742}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000011; Y = 8'b00011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2377,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1742
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111100; Y = 8'b11110111; // Expected: {'Z': -540}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111100; Y = 8'b11110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2378,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110010; Y = 8'b00101000; // Expected: {'Z': 2000}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110010; Y = 8'b00101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2379,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001000; Y = 8'b11100101; // Expected: {'Z': 3240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001000; Y = 8'b11100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2380,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b11110000; // Expected: {'Z': -976}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b11110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2381,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -976
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b01111101; // Expected: {'Z': -7375}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b01111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2382,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7375
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010010; Y = 8'b00100010; // Expected: {'Z': 2788}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010010; Y = 8'b00100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2383,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2788
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000101; Y = 8'b10000010; // Expected: {'Z': -630}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000101; Y = 8'b10000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2384,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -630
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001100; Y = 8'b00010000; // Expected: {'Z': 192}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001100; Y = 8'b00010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2385,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110100; Y = 8'b00010101; // Expected: {'Z': -1596}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110100; Y = 8'b00010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2386,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1596
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011100; Y = 8'b00111000; // Expected: {'Z': 1568}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011100; Y = 8'b00111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2387,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1568
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111000; Y = 8'b00000111; // Expected: {'Z': -56}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111000; Y = 8'b00000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2388,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b11000000; // Expected: {'Z': -1216}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b11000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2389,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110001; Y = 8'b10110011; // Expected: {'Z': 6083}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110001; Y = 8'b10110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2390,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6083
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b01011110; // Expected: {'Z': 5076}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b01011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2391,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5076
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110101; Y = 8'b01100011; // Expected: {'Z': -1089}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110101; Y = 8'b01100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2392,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1089
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b00110000; // Expected: {'Z': -4176}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b00110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2393,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001000; Y = 8'b11100011; // Expected: {'Z': -232}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001000; Y = 8'b11100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2394,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111001; Y = 8'b01100101; // Expected: {'Z': -7171}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111001; Y = 8'b01100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2395,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001010; Y = 8'b00100101; // Expected: {'Z': -4366}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001010; Y = 8'b00100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2396,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4366
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100001; Y = 8'b00110111; // Expected: {'Z': -1705}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100001; Y = 8'b00110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2397,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1705
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b01110010; // Expected: {'Z': 7752}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b01110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2398,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7752
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001010; Y = 8'b01111100; // Expected: {'Z': -6696}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001010; Y = 8'b01111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2399,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6696
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011010; Y = 8'b00011011; // Expected: {'Z': -1026}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011010; Y = 8'b00011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2400,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1026
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010100; Y = 8'b11011010; // Expected: {'Z': 1672}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010100; Y = 8'b11011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2401,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011001; Y = 8'b00111001; // Expected: {'Z': 1425}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011001; Y = 8'b00111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2402,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1425
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b00100110; // Expected: {'Z': 2318}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b00100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2403,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2318
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b00001010; // Expected: {'Z': 1120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b00001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2404,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000001; Y = 8'b00110110; // Expected: {'Z': -6858}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000001; Y = 8'b00110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2405,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6858
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b11101001; // Expected: {'Z': -299}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b11101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2406,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -299
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011110; Y = 8'b11110111; // Expected: {'Z': 306}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011110; Y = 8'b11110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2407,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 306
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111100; Y = 8'b10110000; // Expected: {'Z': -4800}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111100; Y = 8'b10110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2408,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011100; Y = 8'b01001100; // Expected: {'Z': -7600}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011100; Y = 8'b01001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2409,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100010; Y = 8'b01010100; // Expected: {'Z': 2856}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100010; Y = 8'b01010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2410,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010001; Y = 8'b10101001; // Expected: {'Z': 4089}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010001; Y = 8'b10101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2411,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4089
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001100; Y = 8'b10111111; // Expected: {'Z': 3380}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001100; Y = 8'b10111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2412,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3380
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101101; Y = 8'b11010110; // Expected: {'Z': 798}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101101; Y = 8'b11010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2413,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101100; Y = 8'b00110001; // Expected: {'Z': -980}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101100; Y = 8'b00110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2414,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100000; Y = 8'b10101100; // Expected: {'Z': -2688}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100000; Y = 8'b10101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2415,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2688
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110000; Y = 8'b11100100; // Expected: {'Z': 448}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110000; Y = 8'b11100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2416,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 448
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001100; Y = 8'b01111011; // Expected: {'Z': -14268}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001100; Y = 8'b01111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2417,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -14268
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111001; Y = 8'b00111001; // Expected: {'Z': -399}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111001; Y = 8'b00111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2418,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -399
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010111; Y = 8'b00111010; // Expected: {'Z': 1334}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010111; Y = 8'b00111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2419,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1334
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010011; Y = 8'b10110011; // Expected: {'Z': -6391}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010011; Y = 8'b10110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2420,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6391
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010111; Y = 8'b00110001; // Expected: {'Z': -2009}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010111; Y = 8'b00110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2421,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2009
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b10110101; // Expected: {'Z': -4575}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b10110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2422,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4575
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010111; Y = 8'b11001101; // Expected: {'Z': 2091}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010111; Y = 8'b11001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2423,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2091
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b01001111; // Expected: {'Z': 158}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b01001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2424,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 158
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001010; Y = 8'b11011111; // Expected: {'Z': 1782}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001010; Y = 8'b11011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2425,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1782
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010100; Y = 8'b10010110; // Expected: {'Z': -8904}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010100; Y = 8'b10010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2426,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8904
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b01010110; // Expected: {'Z': 5246}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b01010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2427,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111101; Y = 8'b00110010; // Expected: {'Z': 6250}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111101; Y = 8'b00110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2428,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110010; Y = 8'b11010111; // Expected: {'Z': -4674}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110010; Y = 8'b11010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2429,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4674
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b10110001; // Expected: {'Z': 4029}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b10110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2430,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4029
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111110; Y = 8'b10110111; // Expected: {'Z': 146}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111110; Y = 8'b10110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2431,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101001; Y = 8'b10111001; // Expected: {'Z': -2911}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101001; Y = 8'b10111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2432,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2911
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001011; Y = 8'b01000100; // Expected: {'Z': -7956}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001011; Y = 8'b01000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2433,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7956
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b10011111; // Expected: {'Z': -582}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b10011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2434,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -582
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111011; Y = 8'b01011000; // Expected: {'Z': -6072}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111011; Y = 8'b01011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2435,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6072
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000010; Y = 8'b01101100; // Expected: {'Z': -13608}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000010; Y = 8'b01101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2436,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -13608
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000001; Y = 8'b10010011; // Expected: {'Z': 13843}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000001; Y = 8'b10010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2437,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 13843
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101010; Y = 8'b11000001; // Expected: {'Z': 1386}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101010; Y = 8'b11000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2438,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1386
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001101; Y = 8'b10010110; // Expected: {'Z': -8162}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001101; Y = 8'b10010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2439,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011111; Y = 8'b01011100; // Expected: {'Z': 8740}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011111; Y = 8'b01011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2440,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8740
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111010; Y = 8'b00011011; // Expected: {'Z': -162}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111010; Y = 8'b00011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2441,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110011; Y = 8'b11011011; // Expected: {'Z': 481}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110011; Y = 8'b11011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2442,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 481
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b11111100; // Expected: {'Z': 328}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b11111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2443,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 328
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000100; Y = 8'b01100111; // Expected: {'Z': -6180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000100; Y = 8'b01100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2444,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111011; Y = 8'b11010010; // Expected: {'Z': -2714}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111011; Y = 8'b11010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2445,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2714
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111000; Y = 8'b11011001; // Expected: {'Z': 2808}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111000; Y = 8'b11011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2446,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100100; Y = 8'b01100001; // Expected: {'Z': -8924}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100100; Y = 8'b01100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2447,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8924
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001100; Y = 8'b00101101; // Expected: {'Z': 540}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001100; Y = 8'b00101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2448,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000110; Y = 8'b11101100; // Expected: {'Z': 1160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000110; Y = 8'b11101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2449,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001110; Y = 8'b10001100; // Expected: {'Z': 5800}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001110; Y = 8'b10001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2450,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001010; Y = 8'b11000110; // Expected: {'Z': -580}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001010; Y = 8'b11000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2451,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110100; Y = 8'b11111111; // Expected: {'Z': -52}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110100; Y = 8'b11111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2452,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111000; Y = 8'b11110001; // Expected: {'Z': 120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111000; Y = 8'b11110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2453,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110010; Y = 8'b10000011; // Expected: {'Z': 1750}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110010; Y = 8'b10000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2454,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111000; Y = 8'b01110010; // Expected: {'Z': -912}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111000; Y = 8'b01110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2455,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -912
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000001; Y = 8'b01101100; // Expected: {'Z': -6804}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000001; Y = 8'b01101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2456,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6804
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000100; Y = 8'b10011111; // Expected: {'Z': -388}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000100; Y = 8'b10011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2457,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -388
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110001; Y = 8'b01110110; // Expected: {'Z': -1770}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110001; Y = 8'b01110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2458,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1770
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101010; Y = 8'b10001101; // Expected: {'Z': -4830}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101010; Y = 8'b10001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2459,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4830
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001100; Y = 8'b10010011; // Expected: {'Z': 12644}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001100; Y = 8'b10010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2460,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 12644
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100011; Y = 8'b10111011; // Expected: {'Z': 2001}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100011; Y = 8'b10111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2461,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2001
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010000; Y = 8'b00001001; // Expected: {'Z': 144}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010000; Y = 8'b00001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2462,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b01000010; // Expected: {'Z': -3366}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b01000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2463,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3366
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b10001010; // Expected: {'Z': -1534}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b10001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2464,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1534
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100000; Y = 8'b11111001; // Expected: {'Z': 672}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100000; Y = 8'b11111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2465,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110001; Y = 8'b00111101; // Expected: {'Z': -915}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110001; Y = 8'b00111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2466,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -915
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b00011100; // Expected: {'Z': 2884}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b00011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2467,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2884
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000111; Y = 8'b01110110; // Expected: {'Z': 826}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000111; Y = 8'b01110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2468,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 826
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111110; Y = 8'b11000001; // Expected: {'Z': 4158}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111110; Y = 8'b11000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2469,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4158
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100000; Y = 8'b00111000; // Expected: {'Z': 1792}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100000; Y = 8'b00111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2470,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101011; Y = 8'b00111001; // Expected: {'Z': -4845}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101011; Y = 8'b00111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2471,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4845
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011101; Y = 8'b10010001; // Expected: {'Z': 3885}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011101; Y = 8'b10010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2472,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3885
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011000; Y = 8'b11010100; // Expected: {'Z': -1056}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011000; Y = 8'b11010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2473,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1056
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101010; Y = 8'b10011011; // Expected: {'Z': 2222}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101010; Y = 8'b10011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2474,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100110; Y = 8'b10011100; // Expected: {'Z': 2600}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100110; Y = 8'b10011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2475,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100000; Y = 8'b11100010; // Expected: {'Z': 960}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100000; Y = 8'b11100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2476,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111001; Y = 8'b10110100; // Expected: {'Z': 5396}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111001; Y = 8'b10110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2477,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5396
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111001; Y = 8'b01100011; // Expected: {'Z': 5643}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111001; Y = 8'b01100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2478,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5643
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010100; Y = 8'b01100110; // Expected: {'Z': 8568}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010100; Y = 8'b01100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2479,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8568
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000011; Y = 8'b10010000; // Expected: {'Z': -336}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000011; Y = 8'b10010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2480,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -336
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011010; Y = 8'b01011110; // Expected: {'Z': 8460}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011010; Y = 8'b01011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2481,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8460
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010000; Y = 8'b01110101; // Expected: {'Z': -5616}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010000; Y = 8'b01110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2482,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5616
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100111; Y = 8'b00100110; // Expected: {'Z': -3382}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100111; Y = 8'b00100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2483,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3382
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010010; Y = 8'b10101101; // Expected: {'Z': -6806}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010010; Y = 8'b10101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2484,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6806
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101000; Y = 8'b10010100; // Expected: {'Z': 2592}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101000; Y = 8'b10010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2485,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2592
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100011; Y = 8'b01000111; // Expected: {'Z': 2485}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100011; Y = 8'b01000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2486,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2485
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111000; Y = 8'b10111111; // Expected: {'Z': -3640}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111000; Y = 8'b10111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2487,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101001; Y = 8'b11110111; // Expected: {'Z': -369}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101001; Y = 8'b11110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2488,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -369
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010000; Y = 8'b00001101; // Expected: {'Z': -1456}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010000; Y = 8'b00001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2489,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000101; Y = 8'b10101000; // Expected: {'Z': -440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000101; Y = 8'b10101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2490,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101100; Y = 8'b00000111; // Expected: {'Z': -140}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101100; Y = 8'b00000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2491,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001111; Y = 8'b01000110; // Expected: {'Z': -3430}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001111; Y = 8'b01000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2492,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001100; Y = 8'b01100110; // Expected: {'Z': -11832}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001100; Y = 8'b01100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2493,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11832
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100010; Y = 8'b10111010; // Expected: {'Z': 2100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100010; Y = 8'b10111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2494,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110011; Y = 8'b01101000; // Expected: {'Z': -1352}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110011; Y = 8'b01101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2495,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111011; Y = 8'b01001010; // Expected: {'Z': -370}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111011; Y = 8'b01001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2496,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -370
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000000; Y = 8'b11000100; // Expected: {'Z': 3840}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000000; Y = 8'b11000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2497,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001100; Y = 8'b11101010; // Expected: {'Z': 1144}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001100; Y = 8'b11101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2498,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110000; Y = 8'b11001100; // Expected: {'Z': -2496}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110000; Y = 8'b11001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2499,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100000; Y = 8'b10100000; // Expected: {'Z': -3072}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100000; Y = 8'b10100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2500,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3072
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110000; Y = 8'b00101000; // Expected: {'Z': 1920}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110000; Y = 8'b00101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2501,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011010; Y = 8'b00001001; // Expected: {'Z': -918}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011010; Y = 8'b00001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2502,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -918
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b11000010; // Expected: {'Z': -6944}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b11000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2503,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111000; Y = 8'b00111001; // Expected: {'Z': 3192}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111000; Y = 8'b00111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2504,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010011; Y = 8'b00000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010011; Y = 8'b00000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2505,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010000; Y = 8'b01101011; // Expected: {'Z': 1712}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010000; Y = 8'b01101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2506,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1712
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101111; Y = 8'b11010110; // Expected: {'Z': 714}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101111; Y = 8'b11010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2507,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 714
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001101; Y = 8'b10111011; // Expected: {'Z': 7935}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001101; Y = 8'b10111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2508,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7935
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011001; Y = 8'b00010111; // Expected: {'Z': -897}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011001; Y = 8'b00010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2509,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -897
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000100; Y = 8'b00011010; // Expected: {'Z': 104}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000100; Y = 8'b00011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2510,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100100; Y = 8'b00011111; // Expected: {'Z': -2852}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100100; Y = 8'b00011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2511,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2852
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001011; Y = 8'b01101010; // Expected: {'Z': -5618}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001011; Y = 8'b01101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2512,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5618
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010111; Y = 8'b01100111; // Expected: {'Z': -10815}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010111; Y = 8'b01100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2513,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10815
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111011; Y = 8'b00010000; // Expected: {'Z': 944}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111011; Y = 8'b00010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2514,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110011; Y = 8'b01111100; // Expected: {'Z': -9548}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110011; Y = 8'b01111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2515,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9548
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110011; Y = 8'b01100111; // Expected: {'Z': 5253}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110011; Y = 8'b01100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2516,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000110; Y = 8'b01111010; // Expected: {'Z': -14884}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000110; Y = 8'b01111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2517,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -14884
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010100; Y = 8'b01111111; // Expected: {'Z': -13716}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010100; Y = 8'b01111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2518,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -13716
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111101; Y = 8'b11001110; // Expected: {'Z': 150}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111101; Y = 8'b11001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2519,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010100; Y = 8'b10010001; // Expected: {'Z': 11988}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010100; Y = 8'b10010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2520,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11988
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110011; Y = 8'b01011011; // Expected: {'Z': 4641}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110011; Y = 8'b01011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2521,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4641
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b10011011; // Expected: {'Z': -4444}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b10011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2522,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4444
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010001; Y = 8'b01101000; // Expected: {'Z': 8424}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010001; Y = 8'b01101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2523,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8424
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010110; Y = 8'b00111011; // Expected: {'Z': 5074}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010110; Y = 8'b00111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2524,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5074
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110101; Y = 8'b00101010; // Expected: {'Z': -3150}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110101; Y = 8'b00101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2525,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b00100001; // Expected: {'Z': 627}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b00100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2526,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 627
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011001; Y = 8'b11111111; // Expected: {'Z': -89}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011001; Y = 8'b11111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2527,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -89
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b00101011; // Expected: {'Z': -2408}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b00101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2528,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001000; Y = 8'b11111011; // Expected: {'Z': -40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001000; Y = 8'b11111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2529,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011110; Y = 8'b00000111; // Expected: {'Z': -238}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011110; Y = 8'b00000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2530,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111110; Y = 8'b00011000; // Expected: {'Z': 1488}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111110; Y = 8'b00011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2531,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b00010011; // Expected: {'Z': -532}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b00010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2532,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -532
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000111; Y = 8'b00011111; // Expected: {'Z': 2201}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000111; Y = 8'b00011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2533,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000011; Y = 8'b11111110; // Expected: {'Z': -6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000011; Y = 8'b11111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2534,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b11010000; // Expected: {'Z': -288}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b11010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2535,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011011; Y = 8'b01010000; // Expected: {'Z': 2160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011011; Y = 8'b01010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2536,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b11000011; // Expected: {'Z': -915}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b11000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2537,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -915
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b01001001; // Expected: {'Z': -4307}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b01001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2538,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4307
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100010; Y = 8'b01001001; // Expected: {'Z': -6862}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100010; Y = 8'b01001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2539,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6862
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111101; Y = 8'b00010110; // Expected: {'Z': -1474}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111101; Y = 8'b00010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2540,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1474
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101001; Y = 8'b10000010; // Expected: {'Z': -13230}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101001; Y = 8'b10000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2541,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -13230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b00010010; // Expected: {'Z': 522}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b00010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2542,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 522
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011110; Y = 8'b01100111; // Expected: {'Z': 9682}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011110; Y = 8'b01100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2543,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9682
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010100; Y = 8'b00000111; // Expected: {'Z': 140}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010100; Y = 8'b00000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2544,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010100; Y = 8'b00101000; // Expected: {'Z': -4320}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010100; Y = 8'b00101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2545,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b00010001; // Expected: {'Z': 612}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b00010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2546,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110001; Y = 8'b00101110; // Expected: {'Z': 2254}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110001; Y = 8'b00101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2547,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011110; Y = 8'b01110100; // Expected: {'Z': -11368}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011110; Y = 8'b01110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2548,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011011; Y = 8'b01001011; // Expected: {'Z': 6825}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011011; Y = 8'b01001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2549,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6825
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111001; Y = 8'b00010011; // Expected: {'Z': 1083}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111001; Y = 8'b00010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2550,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1083
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b10101010; // Expected: {'Z': -4644}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b10101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2551,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4644
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000110; Y = 8'b10110111; // Expected: {'Z': 8906}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000110; Y = 8'b10110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2552,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8906
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b10010001; // Expected: {'Z': 9657}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b10010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2553,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9657
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000010; Y = 8'b01101110; // Expected: {'Z': -6820}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000010; Y = 8'b01101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2554,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100101; Y = 8'b01110000; // Expected: {'Z': 4144}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100101; Y = 8'b01110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2555,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001010; Y = 8'b00111101; // Expected: {'Z': 610}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001010; Y = 8'b00111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2556,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 610
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011100; Y = 8'b00001111; // Expected: {'Z': 420}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011100; Y = 8'b00001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2557,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001101; Y = 8'b10100010; // Expected: {'Z': -7238}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001101; Y = 8'b10100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2558,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001111; Y = 8'b00111010; // Expected: {'Z': -6554}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001111; Y = 8'b00111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2559,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6554
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b00101101; // Expected: {'Z': -2655}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b00101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2560,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2655
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111001; Y = 8'b10111101; // Expected: {'Z': 469}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111001; Y = 8'b10111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2561,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 469
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000000; Y = 8'b10011100; // Expected: {'Z': 6400}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000000; Y = 8'b10011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2562,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100000; Y = 8'b00111001; // Expected: {'Z': 1824}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100000; Y = 8'b00111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2563,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1824
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001011; Y = 8'b11001010; // Expected: {'Z': 6318}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001011; Y = 8'b11001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2564,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6318
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b01110000; // Expected: {'Z': -7616}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b01110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2565,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7616
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b10011000; // Expected: {'Z': -7072}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b10011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2566,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7072
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001110; Y = 8'b01011101; // Expected: {'Z': 1302}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001110; Y = 8'b01011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2567,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1302
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000110; Y = 8'b11100100; // Expected: {'Z': 3416}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000110; Y = 8'b11100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2568,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000011; Y = 8'b11111010; // Expected: {'Z': 366}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000011; Y = 8'b11111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2569,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 366
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000001; Y = 8'b01111101; // Expected: {'Z': -7875}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000001; Y = 8'b01111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2570,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7875
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001100; Y = 8'b10101010; // Expected: {'Z': 4472}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001100; Y = 8'b10101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2571,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4472
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110000; Y = 8'b11100011; // Expected: {'Z': -1392}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110000; Y = 8'b11100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2572,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101000; Y = 8'b00101001; // Expected: {'Z': 4264}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101000; Y = 8'b00101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2573,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110100; Y = 8'b01010001; // Expected: {'Z': -972}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110100; Y = 8'b01010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2574,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -972
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010101; Y = 8'b10100001; // Expected: {'Z': 10165}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010101; Y = 8'b10100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2575,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b01111011; // Expected: {'Z': -3444}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b01111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2576,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3444
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b11001101; // Expected: {'Z': -459}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b11001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2577,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -459
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b00010010; // Expected: {'Z': 1224}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b00010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2578,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011111; Y = 8'b10110000; // Expected: {'Z': -7600}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011111; Y = 8'b10110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2579,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101001; Y = 8'b11001011; // Expected: {'Z': 1219}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101001; Y = 8'b11001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2580,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1219
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000001; Y = 8'b11111101; // Expected: {'Z': -3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000001; Y = 8'b11111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2581,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000001; Y = 8'b10001010; // Expected: {'Z': -7670}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000001; Y = 8'b10001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2582,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7670
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010011; Y = 8'b01111101; // Expected: {'Z': 10375}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010011; Y = 8'b01111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2583,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10375
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011010; Y = 8'b11001110; // Expected: {'Z': 1900}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011010; Y = 8'b11001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2584,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111110; Y = 8'b11001111; // Expected: {'Z': -3038}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111110; Y = 8'b11001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2585,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3038
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111101; Y = 8'b00000011; // Expected: {'Z': -9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111101; Y = 8'b00000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2586,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b10011010; // Expected: {'Z': -12546}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b10011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2587,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111110; Y = 8'b01111111; // Expected: {'Z': -254}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111110; Y = 8'b01111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2588,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011011; Y = 8'b01010011; // Expected: {'Z': 7553}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011011; Y = 8'b01010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2589,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7553
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010100; Y = 8'b10110111; // Expected: {'Z': 7884}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010100; Y = 8'b10110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2590,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7884
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100011; Y = 8'b11100011; // Expected: {'Z': 841}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100011; Y = 8'b11100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2591,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 841
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101000; Y = 8'b11111000; // Expected: {'Z': 192}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101000; Y = 8'b11111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2592,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010111; Y = 8'b10011110; // Expected: {'Z': -8526}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010111; Y = 8'b10011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2593,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8526
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010010; Y = 8'b00101101; // Expected: {'Z': 3690}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010010; Y = 8'b00101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2594,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3690
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b10001110; // Expected: {'Z': -11742}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b10001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2595,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11742
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010001; Y = 8'b00001001; // Expected: {'Z': 729}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010001; Y = 8'b00001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2596,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 729
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010111; Y = 8'b01100100; // Expected: {'Z': 8700}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010111; Y = 8'b01100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2597,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001110; Y = 8'b01110100; // Expected: {'Z': -13224}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001110; Y = 8'b01110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2598,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -13224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101000; Y = 8'b00000001; // Expected: {'Z': -88}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101000; Y = 8'b00000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2599,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100001; Y = 8'b11011001; // Expected: {'Z': 1209}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100001; Y = 8'b11011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2600,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b10111100; // Expected: {'Z': -1292}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b10111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2601,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1292
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111110; Y = 8'b10100010; // Expected: {'Z': -5828}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111110; Y = 8'b10100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2602,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101110; Y = 8'b00111100; // Expected: {'Z': 2760}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101110; Y = 8'b00111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2603,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100101; Y = 8'b10111100; // Expected: {'Z': 1836}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100101; Y = 8'b10111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2604,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1836
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010110; Y = 8'b01110001; // Expected: {'Z': -4746}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010110; Y = 8'b01110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2605,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4746
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011110; Y = 8'b00110010; // Expected: {'Z': 4700}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011110; Y = 8'b00110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2606,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b00001110; // Expected: {'Z': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b00001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2607,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010010; Y = 8'b10011101; // Expected: {'Z': -8118}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010010; Y = 8'b10011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2608,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b10010101; // Expected: {'Z': -2033}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b10010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2609,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2033
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b00111010; // Expected: {'Z': 3538}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b00111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2610,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3538
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000000; Y = 8'b00101010; // Expected: {'Z': -5376}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000000; Y = 8'b00101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2611,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5376
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b11110101; // Expected: {'Z': -242}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b11110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2612,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010001; Y = 8'b10110111; // Expected: {'Z': -1241}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010001; Y = 8'b10110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2613,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001100; Y = 8'b00110111; // Expected: {'Z': 660}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001100; Y = 8'b00110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2614,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110011; Y = 8'b00101101; // Expected: {'Z': 5175}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110011; Y = 8'b00101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2615,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000000; Y = 8'b00101100; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000000; Y = 8'b00101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2616,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000100; Y = 8'b00001000; // Expected: {'Z': -480}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000100; Y = 8'b00001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2617,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011100; Y = 8'b01011110; // Expected: {'Z': -9400}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011100; Y = 8'b01011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2618,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111000; Y = 8'b11010001; // Expected: {'Z': 3384}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111000; Y = 8'b11010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2619,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3384
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110010; Y = 8'b11000001; // Expected: {'Z': -3150}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110010; Y = 8'b11000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2620,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101100; Y = 8'b00101100; // Expected: {'Z': -880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101100; Y = 8'b00101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2621,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101100; Y = 8'b00110011; // Expected: {'Z': -1020}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101100; Y = 8'b00110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2622,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1020
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111111; Y = 8'b00111011; // Expected: {'Z': -59}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111111; Y = 8'b00111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2623,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b10111010; // Expected: {'Z': -4760}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b10111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2624,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b11100110; // Expected: {'Z': -52}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b11100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2625,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111011; Y = 8'b00101010; // Expected: {'Z': -210}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111011; Y = 8'b00101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2626,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110101; Y = 8'b01110000; // Expected: {'Z': 5936}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110101; Y = 8'b01110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2627,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5936
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010100; Y = 8'b01000111; // Expected: {'Z': 5964}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010100; Y = 8'b01000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2628,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5964
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001001; Y = 8'b00000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001001; Y = 8'b00000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2629,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100001; Y = 8'b10111111; // Expected: {'Z': 6175}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100001; Y = 8'b10111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2630,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101111; Y = 8'b10000100; // Expected: {'Z': 2108}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101111; Y = 8'b10000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2631,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b01100011; // Expected: {'Z': -5544}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b01100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2632,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5544
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000000; Y = 8'b01110100; // Expected: {'Z': 7424}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000000; Y = 8'b01110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2633,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7424
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b10100101; // Expected: {'Z': 10101}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b10100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2634,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101010; Y = 8'b10010001; // Expected: {'Z': 9546}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101010; Y = 8'b10010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2635,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010001; Y = 8'b01101000; // Expected: {'Z': -4888}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010001; Y = 8'b01101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2636,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010010; Y = 8'b10101100; // Expected: {'Z': 3864}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010010; Y = 8'b10101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2637,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3864
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101111; Y = 8'b10110110; // Expected: {'Z': 1258}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101111; Y = 8'b10110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2638,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1258
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001110; Y = 8'b10110011; // Expected: {'Z': -6006}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001110; Y = 8'b10110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2639,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6006
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b00001100; // Expected: {'Z': -672}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b00001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2640,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b11000000; // Expected: {'Z': 3584}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b11000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2641,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3584
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100110; Y = 8'b01000100; // Expected: {'Z': 6936}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100110; Y = 8'b01000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2642,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6936
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010101; Y = 8'b11111110; // Expected: {'Z': -170}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010101; Y = 8'b11111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2643,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110101; Y = 8'b00110110; // Expected: {'Z': 2862}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110101; Y = 8'b00110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2644,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2862
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011110; Y = 8'b11111010; // Expected: {'Z': -564}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011110; Y = 8'b11111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2645,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -564
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000110; Y = 8'b00110010; // Expected: {'Z': 3500}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000110; Y = 8'b00110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2646,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110000; Y = 8'b00110011; // Expected: {'Z': 2448}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110000; Y = 8'b00110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2647,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2448
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110001; Y = 8'b10100100; // Expected: {'Z': 7268}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110001; Y = 8'b10100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2648,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7268
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011110; Y = 8'b10111111; // Expected: {'Z': 6370}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011110; Y = 8'b10111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2649,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6370
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110100; Y = 8'b00001111; // Expected: {'Z': -180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110100; Y = 8'b00001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2650,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011010; Y = 8'b11010111; // Expected: {'Z': -1066}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011010; Y = 8'b11010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2651,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1066
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101101; Y = 8'b01011010; // Expected: {'Z': 4050}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101101; Y = 8'b01011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2652,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000000; Y = 8'b01101000; // Expected: {'Z': -13312}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000000; Y = 8'b01101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2653,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -13312
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001110; Y = 8'b11011100; // Expected: {'Z': 4104}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001110; Y = 8'b11011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2654,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100111; Y = 8'b01111100; // Expected: {'Z': -11036}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100111; Y = 8'b01111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2655,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11036
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011100; Y = 8'b10001010; // Expected: {'Z': 4248}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011100; Y = 8'b10001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2656,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010111; Y = 8'b11100011; // Expected: {'Z': 3045}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010111; Y = 8'b11100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2657,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3045
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010111; Y = 8'b11001100; // Expected: {'Z': 5460}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010111; Y = 8'b11001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2658,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5460
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011011; Y = 8'b00110111; // Expected: {'Z': -5555}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011011; Y = 8'b00110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2659,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5555
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001001; Y = 8'b10100010; // Expected: {'Z': 5170}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001001; Y = 8'b10100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2660,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000001; Y = 8'b00110110; // Expected: {'Z': -6858}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000001; Y = 8'b00110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2661,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6858
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000010; Y = 8'b10011011; // Expected: {'Z': 12726}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000010; Y = 8'b10011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2662,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 12726
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b01101101; // Expected: {'Z': -7412}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b01101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2663,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7412
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110100; Y = 8'b11101010; // Expected: {'Z': 264}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110100; Y = 8'b11101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2664,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111100; Y = 8'b00110111; // Expected: {'Z': 3300}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111100; Y = 8'b00110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2665,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000100; Y = 8'b01011100; // Expected: {'Z': 368}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000100; Y = 8'b01011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2666,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010111; Y = 8'b11110010; // Expected: {'Z': 1470}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010111; Y = 8'b11110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2667,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1470
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110010; Y = 8'b01101100; // Expected: {'Z': 12312}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110010; Y = 8'b01101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2668,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 12312
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100010; Y = 8'b10110011; // Expected: {'Z': -2618}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100010; Y = 8'b10110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2669,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2618
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101001; Y = 8'b10001100; // Expected: {'Z': -12180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101001; Y = 8'b10001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2670,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100010; Y = 8'b01010111; // Expected: {'Z': 2958}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100010; Y = 8'b01010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2671,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2958
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110101; Y = 8'b11010110; // Expected: {'Z': -4914}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110101; Y = 8'b11010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2672,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4914
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100011; Y = 8'b10011100; // Expected: {'Z': 9300}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100011; Y = 8'b10011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2673,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010000; Y = 8'b00010100; // Expected: {'Z': 320}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010000; Y = 8'b00010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2674,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111110; Y = 8'b01111100; // Expected: {'Z': -248}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111110; Y = 8'b01111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2675,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100110; Y = 8'b10101111; // Expected: {'Z': -8262}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100110; Y = 8'b10101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2676,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8262
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110101; Y = 8'b00010100; // Expected: {'Z': 2340}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110101; Y = 8'b00010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2677,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101100; Y = 8'b10110100; // Expected: {'Z': 1520}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101100; Y = 8'b10110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2678,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100011; Y = 8'b01010000; // Expected: {'Z': 2800}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100011; Y = 8'b01010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2679,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000110; Y = 8'b01101111; // Expected: {'Z': 7770}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000110; Y = 8'b01101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2680,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7770
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111010; Y = 8'b10111110; // Expected: {'Z': -8052}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111010; Y = 8'b10111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2681,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8052
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001111; Y = 8'b01110011; // Expected: {'Z': 9085}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001111; Y = 8'b01110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2682,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9085
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111011; Y = 8'b11011101; // Expected: {'Z': -2065}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111011; Y = 8'b11011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2683,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2065
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100001; Y = 8'b11000110; // Expected: {'Z': -1914}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100001; Y = 8'b11000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2684,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1914
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000011; Y = 8'b11101101; // Expected: {'Z': 1159}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000011; Y = 8'b11101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2685,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011111; Y = 8'b11010101; // Expected: {'Z': -4085}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011111; Y = 8'b11010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2686,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4085
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010101; Y = 8'b00111101; // Expected: {'Z': -6527}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010101; Y = 8'b00111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2687,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6527
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100111; Y = 8'b01001110; // Expected: {'Z': -6942}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100111; Y = 8'b01001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2688,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6942
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b10111100; // Expected: {'Z': 5712}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b10111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2689,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5712
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110000; Y = 8'b11010101; // Expected: {'Z': -2064}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110000; Y = 8'b11010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2690,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2064
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b00001010; // Expected: {'Z': 130}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b00001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2691,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111010; Y = 8'b11000010; // Expected: {'Z': 372}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111010; Y = 8'b11000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2692,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 372
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b10000011; // Expected: {'Z': -9250}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b10000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2693,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010111; Y = 8'b01100000; // Expected: {'Z': 2208}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010111; Y = 8'b01100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2694,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001000; Y = 8'b00100010; // Expected: {'Z': -4080}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001000; Y = 8'b00100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2695,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010100; Y = 8'b11011000; // Expected: {'Z': 4320}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010100; Y = 8'b11011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2696,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b00110000; // Expected: {'Z': -2448}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b00110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2697,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2448
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b01000011; // Expected: {'Z': -4556}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b01000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2698,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4556
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b01101010; // Expected: {'Z': 4134}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b01101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2699,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101011; Y = 8'b01000010; // Expected: {'Z': -5610}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101011; Y = 8'b01000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2700,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5610
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101111; Y = 8'b01111000; // Expected: {'Z': -2040}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101111; Y = 8'b01111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2701,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001011; Y = 8'b00110011; // Expected: {'Z': 3825}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001011; Y = 8'b00110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2702,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3825
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100101; Y = 8'b11001011; // Expected: {'Z': -5353}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100101; Y = 8'b11001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2703,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5353
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110110; Y = 8'b11100001; // Expected: {'Z': -3658}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110110; Y = 8'b11100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2704,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3658
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101000; Y = 8'b10111100; // Expected: {'Z': 1632}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101000; Y = 8'b10111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2705,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1632
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000000; Y = 8'b01111000; // Expected: {'Z': -15360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000000; Y = 8'b01111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2706,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -15360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101010; Y = 8'b01001111; // Expected: {'Z': -6794}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101010; Y = 8'b01001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2707,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6794
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010101; Y = 8'b10110111; // Expected: {'Z': -6205}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010101; Y = 8'b10110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2708,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101011; Y = 8'b10001010; // Expected: {'Z': -5074}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101011; Y = 8'b10001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2709,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5074
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011001; Y = 8'b00010010; // Expected: {'Z': 450}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011001; Y = 8'b00010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2710,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011100; Y = 8'b10101011; // Expected: {'Z': 8500}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011100; Y = 8'b10101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2711,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111011; Y = 8'b01111110; // Expected: {'Z': 7434}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111011; Y = 8'b01111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2712,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7434
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b00110010; // Expected: {'Z': 750}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b00110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2713,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000001; Y = 8'b00000111; // Expected: {'Z': -441}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000001; Y = 8'b00000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2714,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -441
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001001; Y = 8'b01101101; // Expected: {'Z': -5995}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001001; Y = 8'b01101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2715,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5995
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110010; Y = 8'b10000010; // Expected: {'Z': -6300}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110010; Y = 8'b10000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2716,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b10000010; // Expected: {'Z': -9072}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b10000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2717,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9072
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011111; Y = 8'b00101101; // Expected: {'Z': -4365}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011111; Y = 8'b00101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2718,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4365
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010010; Y = 8'b10110100; // Expected: {'Z': -1368}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010010; Y = 8'b10110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2719,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010100; Y = 8'b10001001; // Expected: {'Z': 12852}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010100; Y = 8'b10001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2720,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 12852
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111111; Y = 8'b10010100; // Expected: {'Z': -6804}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111111; Y = 8'b10010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2721,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6804
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111111; Y = 8'b11110110; // Expected: {'Z': 650}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111111; Y = 8'b11110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2722,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101101; Y = 8'b10001100; // Expected: {'Z': -5220}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101101; Y = 8'b10001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2723,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b00110001; // Expected: {'Z': 931}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b00110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2724,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 931
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b01100000; // Expected: {'Z': 1824}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b01100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2725,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1824
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000000; Y = 8'b01011010; // Expected: {'Z': -5760}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000000; Y = 8'b01011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2726,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b11101111; // Expected: {'Z': 1428}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b11101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2727,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1428
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111111; Y = 8'b00010011; // Expected: {'Z': -1235}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111111; Y = 8'b00010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2728,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1235
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b10001000; // Expected: {'Z': 7080}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b10001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2729,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011100; Y = 8'b11010100; // Expected: {'Z': -1232}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011100; Y = 8'b11010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2730,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010001; Y = 8'b10011101; // Expected: {'Z': -1683}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010001; Y = 8'b10011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2731,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1683
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b10001100; // Expected: {'Z': -11948}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b10001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2732,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11948
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b11011000; // Expected: {'Z': 2240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b11011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2733,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100000; Y = 8'b11000010; // Expected: {'Z': 5952}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100000; Y = 8'b11000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2734,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5952
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b01101101; // Expected: {'Z': -6431}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b01101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2735,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6431
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111010; Y = 8'b10011110; // Expected: {'Z': 588}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111010; Y = 8'b10011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2736,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 588
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101101; Y = 8'b10000011; // Expected: {'Z': -13625}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101101; Y = 8'b10000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2737,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -13625
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000011; Y = 8'b11001000; // Expected: {'Z': -3752}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000011; Y = 8'b11001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2738,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3752
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011000; Y = 8'b01100101; // Expected: {'Z': -10504}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011000; Y = 8'b01100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2739,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b01111001; // Expected: {'Z': -9922}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b01111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2740,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9922
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001010; Y = 8'b00110111; // Expected: {'Z': -6490}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001010; Y = 8'b00110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2741,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6490
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011111; Y = 8'b10001111; // Expected: {'Z': 3729}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011111; Y = 8'b10001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2742,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3729
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111110; Y = 8'b11111111; // Expected: {'Z': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111110; Y = 8'b11111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2743,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010000; Y = 8'b01010101; // Expected: {'Z': 1360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010000; Y = 8'b01010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2744,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110001; Y = 8'b00011111; // Expected: {'Z': -2449}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110001; Y = 8'b00011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2745,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2449
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101111; Y = 8'b01011101; // Expected: {'Z': -7533}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101111; Y = 8'b01011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2746,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7533
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011010; Y = 8'b00001111; // Expected: {'Z': 1350}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011010; Y = 8'b00001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2747,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101111; Y = 8'b00010010; // Expected: {'Z': -1458}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101111; Y = 8'b00010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2748,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1458
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001110; Y = 8'b01001000; // Expected: {'Z': 1008}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001110; Y = 8'b01001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2749,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000000; Y = 8'b10011001; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000000; Y = 8'b10011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2750,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110000; Y = 8'b00011101; // Expected: {'Z': -464}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110000; Y = 8'b00011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2751,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111001; Y = 8'b11110010; // Expected: {'Z': 98}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111001; Y = 8'b11110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2752,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111100; Y = 8'b11110010; // Expected: {'Z': -840}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111100; Y = 8'b11110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2753,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111111; Y = 8'b10101111; // Expected: {'Z': 81}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111111; Y = 8'b10101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2754,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010010; Y = 8'b10001001; // Expected: {'Z': -9758}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010010; Y = 8'b10001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2755,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9758
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b01111001; // Expected: {'Z': -3388}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b01111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2756,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3388
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010010; Y = 8'b10110000; // Expected: {'Z': -1440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010010; Y = 8'b10110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2757,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001101; Y = 8'b11011101; // Expected: {'Z': 4025}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001101; Y = 8'b11011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2758,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4025
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110101; Y = 8'b10010010; // Expected: {'Z': 1210}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110101; Y = 8'b10010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2759,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100101; Y = 8'b01010110; // Expected: {'Z': -2322}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100101; Y = 8'b01010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2760,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2322
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110100; Y = 8'b10111111; // Expected: {'Z': 780}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110100; Y = 8'b10111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2761,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011011; Y = 8'b11010111; // Expected: {'Z': 1517}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011011; Y = 8'b11010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2762,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1517
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b10110110; // Expected: {'Z': -3478}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b10110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2763,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3478
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010010; Y = 8'b10100011; // Expected: {'Z': 10230}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010010; Y = 8'b10100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2764,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100100; Y = 8'b00101101; // Expected: {'Z': -4140}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100100; Y = 8'b00101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2765,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110111; Y = 8'b10111100; // Expected: {'Z': -8092}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110111; Y = 8'b10111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2766,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8092
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b11000011; // Expected: {'Z': -915}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b11000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2767,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -915
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110001; Y = 8'b10111100; // Expected: {'Z': -3332}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110001; Y = 8'b10111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2768,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3332
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001010; Y = 8'b11110100; // Expected: {'Z': 648}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001010; Y = 8'b11110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2769,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000100; Y = 8'b10111101; // Expected: {'Z': -268}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000100; Y = 8'b10111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2770,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -268
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100000; Y = 8'b00110100; // Expected: {'Z': -4992}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100000; Y = 8'b00110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2771,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4992
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011100; Y = 8'b11000000; // Expected: {'Z': -5888}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011100; Y = 8'b11000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2772,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011011; Y = 8'b10000001; // Expected: {'Z': 12827}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011011; Y = 8'b10000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2773,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 12827
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110110; Y = 8'b10100010; // Expected: {'Z': 6956}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110110; Y = 8'b10100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2774,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6956
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100011; Y = 8'b11000010; // Expected: {'Z': -6138}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100011; Y = 8'b11000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2775,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b00000010; // Expected: {'Z': 88}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b00000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2776,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100101; Y = 8'b10111101; // Expected: {'Z': 1809}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100101; Y = 8'b10111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2777,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1809
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110000; Y = 8'b01101011; // Expected: {'Z': -8560}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110000; Y = 8'b01101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2778,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011100; Y = 8'b10110100; // Expected: {'Z': 7600}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011100; Y = 8'b10110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2779,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101001; Y = 8'b00011011; // Expected: {'Z': 1107}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101001; Y = 8'b00011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2780,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b01010111; // Expected: {'Z': 2523}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b01010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2781,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2523
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011101; Y = 8'b11010101; // Expected: {'Z': 4257}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011101; Y = 8'b11010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2782,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4257
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000011; Y = 8'b00000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000011; Y = 8'b00000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2783,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101000; Y = 8'b01010000; // Expected: {'Z': 8320}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101000; Y = 8'b01010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2784,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b01111101; // Expected: {'Z': 9000}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b01111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2785,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101000; Y = 8'b00101111; // Expected: {'Z': -1128}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101000; Y = 8'b00101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2786,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b11110100; // Expected: {'Z': -648}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b11110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2787,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111011; Y = 8'b10110011; // Expected: {'Z': 5313}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111011; Y = 8'b10110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2788,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5313
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b00110110; // Expected: {'Z': -3186}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b00110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2789,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010111; Y = 8'b01111000; // Expected: {'Z': 10440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010111; Y = 8'b01111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2790,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001001; Y = 8'b01101101; // Expected: {'Z': -12971}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001001; Y = 8'b01101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2791,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12971
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b01111100; // Expected: {'Z': 4464}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b01111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2792,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011110; Y = 8'b10111011; // Expected: {'Z': 2346}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011110; Y = 8'b10111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2793,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2346
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110111; Y = 8'b00110101; // Expected: {'Z': 6307}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110111; Y = 8'b00110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2794,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6307
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001111; Y = 8'b10010111; // Expected: {'Z': 5145}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001111; Y = 8'b10010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2795,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010100; Y = 8'b01101101; // Expected: {'Z': -11772}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010100; Y = 8'b01101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2796,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -11772
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001000; Y = 8'b11110111; // Expected: {'Z': -72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001000; Y = 8'b11110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2797,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010011; Y = 8'b00110010; // Expected: {'Z': 4150}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010011; Y = 8'b00110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2798,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011101; Y = 8'b01001100; // Expected: {'Z': -2660}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011101; Y = 8'b01001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2799,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000011; Y = 8'b10101110; // Expected: {'Z': -246}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000011; Y = 8'b10101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2800,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011101; Y = 8'b10011101; // Expected: {'Z': 9801}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011101; Y = 8'b10011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2801,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9801
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011000; Y = 8'b10101010; // Expected: {'Z': 3440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011000; Y = 8'b10101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2802,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110001; Y = 8'b00010100; // Expected: {'Z': 2260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110001; Y = 8'b00010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2803,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101000; Y = 8'b11011101; // Expected: {'Z': -3640}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101000; Y = 8'b11011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2804,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100010; Y = 8'b01110111; // Expected: {'Z': 4046}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100010; Y = 8'b01110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2805,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4046
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111010; Y = 8'b10000011; // Expected: {'Z': 750}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111010; Y = 8'b10000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2806,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b10111000; // Expected: {'Z': 6264}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b10111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2807,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b00010011; // Expected: {'Z': -1596}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b00010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2808,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1596
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100101; Y = 8'b10010100; // Expected: {'Z': -10908}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100101; Y = 8'b10010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2809,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10908
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001010; Y = 8'b11100100; // Expected: {'Z': 3304}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001010; Y = 8'b11100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2810,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3304
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b00101100; // Expected: {'Z': -3696}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b00101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2811,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3696
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b01100011; // Expected: {'Z': 3564}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b01100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2812,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3564
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001111; Y = 8'b01111001; // Expected: {'Z': 9559}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001111; Y = 8'b01111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2813,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9559
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100110; Y = 8'b11100001; // Expected: {'Z': 2790}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100110; Y = 8'b11100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2814,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2790
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001000; Y = 8'b01000110; // Expected: {'Z': 560}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001000; Y = 8'b01000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2815,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001001; Y = 8'b10010011; // Expected: {'Z': -7957}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001001; Y = 8'b10010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2816,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7957
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010101; Y = 8'b01100111; // Expected: {'Z': -4429}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010101; Y = 8'b01100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2817,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4429
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100010; Y = 8'b11000110; // Expected: {'Z': -5684}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100010; Y = 8'b11000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2818,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5684
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001110; Y = 8'b00111000; // Expected: {'Z': 784}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001110; Y = 8'b00111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2819,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011111; Y = 8'b10111100; // Expected: {'Z': -2108}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011111; Y = 8'b10111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2820,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b11111001; // Expected: {'Z': -476}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b11111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2821,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -476
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010010; Y = 8'b10011111; // Expected: {'Z': -1746}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010010; Y = 8'b10011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2822,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1746
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101010; Y = 8'b00001111; // Expected: {'Z': -330}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101010; Y = 8'b00001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2823,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -330
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000000; Y = 8'b11000001; // Expected: {'Z': -4032}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000000; Y = 8'b11000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2824,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4032
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100010; Y = 8'b01000011; // Expected: {'Z': -2010}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100010; Y = 8'b01000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2825,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2010
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000001; Y = 8'b11011010; // Expected: {'Z': -2470}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000001; Y = 8'b11011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2826,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2470
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b11011110; // Expected: {'Z': 2856}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b11011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2827,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b11110101; // Expected: {'Z': -66}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b11110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2828,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111100; Y = 8'b11101100; // Expected: {'Z': -2480}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111100; Y = 8'b11101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2829,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001011; Y = 8'b01111001; // Expected: {'Z': 9075}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001011; Y = 8'b01111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2830,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9075
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b11111110; // Expected: {'Z': -122}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b11111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2831,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100101; Y = 8'b11010010; // Expected: {'Z': 1242}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100101; Y = 8'b11010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2832,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100000; Y = 8'b00000110; // Expected: {'Z': 192}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100000; Y = 8'b00000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2833,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011110; Y = 8'b11010000; // Expected: {'Z': 4704}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011110; Y = 8'b11010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2834,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4704
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011000; Y = 8'b10100011; // Expected: {'Z': 3720}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011000; Y = 8'b10100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2835,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011100; Y = 8'b00001101; // Expected: {'Z': -468}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011100; Y = 8'b00001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2836,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -468
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110011; Y = 8'b10011011; // Expected: {'Z': -5151}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110011; Y = 8'b10011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2837,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5151
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100111; Y = 8'b11000100; // Expected: {'Z': 1500}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100111; Y = 8'b11000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2838,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100100; Y = 8'b00100000; // Expected: {'Z': -2944}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100100; Y = 8'b00100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2839,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010111; Y = 8'b10100100; // Expected: {'Z': 3772}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010111; Y = 8'b10100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2840,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3772
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110110; Y = 8'b11001001; // Expected: {'Z': 4070}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110110; Y = 8'b11001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2841,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4070
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011101; Y = 8'b11010001; // Expected: {'Z': 4653}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011101; Y = 8'b11010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2842,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4653
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101010; Y = 8'b11110011; // Expected: {'Z': 1118}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101010; Y = 8'b11110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2843,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110010; Y = 8'b01011110; // Expected: {'Z': -1316}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110010; Y = 8'b01011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2844,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1316
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100011; Y = 8'b00000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100011; Y = 8'b00000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2845,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100100; Y = 8'b00100000; // Expected: {'Z': 3200}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100100; Y = 8'b00100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2846,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b11000010; // Expected: {'Z': -3348}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b11000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2847,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3348
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101101; Y = 8'b01011001; // Expected: {'Z': -7387}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101101; Y = 8'b01011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2848,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7387
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100000; Y = 8'b00111000; // Expected: {'Z': -5376}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100000; Y = 8'b00111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2849,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5376
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101001; Y = 8'b11101011; // Expected: {'Z': -2205}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101001; Y = 8'b11101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2850,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100011; Y = 8'b10001111; // Expected: {'Z': 3277}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100011; Y = 8'b10001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2851,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3277
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110101; Y = 8'b01000100; // Expected: {'Z': -748}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110101; Y = 8'b01000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2852,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -748
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000001; Y = 8'b11100100; // Expected: {'Z': -1820}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000001; Y = 8'b11100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2853,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b11111100; // Expected: {'Z': -448}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b11111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2854,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -448
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111011; Y = 8'b00111001; // Expected: {'Z': 3363}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111011; Y = 8'b00111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2855,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3363
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001110; Y = 8'b01001110; // Expected: {'Z': -3900}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001110; Y = 8'b01001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2856,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011101; Y = 8'b01111101; // Expected: {'Z': -12375}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011101; Y = 8'b01111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2857,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12375
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111000; Y = 8'b00101010; // Expected: {'Z': -336}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111000; Y = 8'b00101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2858,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -336
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000101; Y = 8'b01010111; // Expected: {'Z': -10701}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000101; Y = 8'b01010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2859,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10701
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010110; Y = 8'b10100111; // Expected: {'Z': 3738}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010110; Y = 8'b10100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2860,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3738
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b10100001; // Expected: {'Z': -3705}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b10100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2861,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3705
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110000; Y = 8'b00111101; // Expected: {'Z': -4880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110000; Y = 8'b00111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2862,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011100; Y = 8'b10000010; // Expected: {'Z': 4536}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011100; Y = 8'b10000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2863,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4536
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010011; Y = 8'b01110110; // Expected: {'Z': -5310}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010011; Y = 8'b01110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2864,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5310
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111001; Y = 8'b10011111; // Expected: {'Z': 6887}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111001; Y = 8'b10011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2865,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6887
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001111; Y = 8'b11001011; // Expected: {'Z': -4187}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001111; Y = 8'b11001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2866,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110000; Y = 8'b00110110; // Expected: {'Z': -864}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110000; Y = 8'b00110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2867,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -864
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000111; Y = 8'b01010010; // Expected: {'Z': 5822}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000111; Y = 8'b01010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2868,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5822
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111010; Y = 8'b10110011; // Expected: {'Z': 462}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111010; Y = 8'b10110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2869,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011010; Y = 8'b10011010; // Expected: {'Z': 3876}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011010; Y = 8'b10011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2870,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3876
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101010; Y = 8'b10001001; // Expected: {'Z': -12614}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101010; Y = 8'b10001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2871,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12614
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001000; Y = 8'b10101110; // Expected: {'Z': 9840}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001000; Y = 8'b10101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2872,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011111; Y = 8'b01010010; // Expected: {'Z': -7954}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011111; Y = 8'b01010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2873,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7954
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b11001100; // Expected: {'Z': -676}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b11001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2874,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -676
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011101; Y = 8'b10010101; // Expected: {'Z': 3745}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011101; Y = 8'b10010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2875,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3745
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010101; Y = 8'b00001100; // Expected: {'Z': 1020}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010101; Y = 8'b00001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2876,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1020
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100101; Y = 8'b10110100; // Expected: {'Z': -7676}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100101; Y = 8'b10110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2877,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7676
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000000; Y = 8'b10110110; // Expected: {'Z': 9472}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000000; Y = 8'b10110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2878,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9472
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000001; Y = 8'b11010010; // Expected: {'Z': 5842}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000001; Y = 8'b11010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2879,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5842
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110000; Y = 8'b11011000; // Expected: {'Z': 640}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110000; Y = 8'b11011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2880,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010100; Y = 8'b10100010; // Expected: {'Z': 4136}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010100; Y = 8'b10100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2881,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b10101111; // Expected: {'Z': -9072}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b10101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2882,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9072
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000010; Y = 8'b00011010; // Expected: {'Z': -3276}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000010; Y = 8'b00011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2883,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3276
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111101; Y = 8'b00000101; // Expected: {'Z': 625}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111101; Y = 8'b00000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2884,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 625
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111001; Y = 8'b11100000; // Expected: {'Z': -3872}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111001; Y = 8'b11100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2885,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3872
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101000; Y = 8'b00001111; // Expected: {'Z': -360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101000; Y = 8'b00001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2886,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101011; Y = 8'b10001110; // Expected: {'Z': 2394}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101011; Y = 8'b10001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2887,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2394
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000011; Y = 8'b11110111; // Expected: {'Z': -603}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000011; Y = 8'b11110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2888,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -603
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001110; Y = 8'b00101111; // Expected: {'Z': 658}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001110; Y = 8'b00101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2889,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 658
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b00111001; // Expected: {'Z': 6384}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b00111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2890,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6384
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001101; Y = 8'b11111110; // Expected: {'Z': -154}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001101; Y = 8'b11111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2891,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110000; Y = 8'b01110110; // Expected: {'Z': 5664}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110000; Y = 8'b01110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2892,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5664
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000011; Y = 8'b11111011; // Expected: {'Z': -335}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000011; Y = 8'b11111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2893,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -335
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011011; Y = 8'b10111111; // Expected: {'Z': 2405}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011011; Y = 8'b10111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2894,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2405
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110001; Y = 8'b10010000; // Expected: {'Z': -5488}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110001; Y = 8'b10010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2895,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100100; Y = 8'b10001110; // Expected: {'Z': 10488}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100100; Y = 8'b10001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2896,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000111; Y = 8'b00111110; // Expected: {'Z': -7502}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000111; Y = 8'b00111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2897,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7502
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001100; Y = 8'b11101110; // Expected: {'Z': -216}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001100; Y = 8'b11101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2898,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101101; Y = 8'b00000111; // Expected: {'Z': 763}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101101; Y = 8'b00000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2899,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 763
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100101; Y = 8'b10001111; // Expected: {'Z': -4181}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100101; Y = 8'b10001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2900,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010011; Y = 8'b00111111; // Expected: {'Z': -2835}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010011; Y = 8'b00111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2901,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2835
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111000; Y = 8'b01110001; // Expected: {'Z': 13560}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111000; Y = 8'b01110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2902,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 13560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011110; Y = 8'b10110101; // Expected: {'Z': 7350}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011110; Y = 8'b10110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2903,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011100; Y = 8'b10001111; // Expected: {'Z': -10396}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011100; Y = 8'b10001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2904,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10396
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011000; Y = 8'b10110100; // Expected: {'Z': 3040}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011000; Y = 8'b10110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2905,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b10110001; // Expected: {'Z': -1027}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b10110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2906,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1027
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010110; Y = 8'b10101101; // Expected: {'Z': 8798}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010110; Y = 8'b10101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2907,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100001; Y = 8'b00001111; // Expected: {'Z': 495}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100001; Y = 8'b00001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2908,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 495
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100101; Y = 8'b10101100; // Expected: {'Z': -3108}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100101; Y = 8'b10101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2909,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010001; Y = 8'b11011000; // Expected: {'Z': 1880}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010001; Y = 8'b11011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2910,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001111; Y = 8'b10000001; // Expected: {'Z': 6223}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001111; Y = 8'b10000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2911,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6223
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011111; Y = 8'b11001011; // Expected: {'Z': 5141}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011111; Y = 8'b11001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2912,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100111; Y = 8'b10110111; // Expected: {'Z': 1825}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100111; Y = 8'b10110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2913,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1825
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111011; Y = 8'b11010100; // Expected: {'Z': 220}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111011; Y = 8'b11010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2914,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011111; Y = 8'b11010010; // Expected: {'Z': 1518}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011111; Y = 8'b11010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2915,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1518
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100101; Y = 8'b00110001; // Expected: {'Z': 1813}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100101; Y = 8'b00110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2916,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1813
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110101; Y = 8'b01000101; // Expected: {'Z': 8073}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110101; Y = 8'b01000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2917,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8073
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011001; Y = 8'b11110101; // Expected: {'Z': -979}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011001; Y = 8'b11110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2918,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -979
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110010; Y = 8'b01001100; // Expected: {'Z': -5928}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110010; Y = 8'b01001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2919,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5928
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010100; Y = 8'b10110010; // Expected: {'Z': 3432}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010100; Y = 8'b10110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2920,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011000; Y = 8'b00100001; // Expected: {'Z': 792}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011000; Y = 8'b00100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2921,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101000; Y = 8'b01100101; // Expected: {'Z': 4040}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101000; Y = 8'b01100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2922,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000111; Y = 8'b10011010; // Expected: {'Z': 5814}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000111; Y = 8'b10011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2923,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5814
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b01101001; // Expected: {'Z': 7560}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b01101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2924,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010110; Y = 8'b11110111; // Expected: {'Z': -774}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010110; Y = 8'b11110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2925,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -774
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100000; Y = 8'b11110001; // Expected: {'Z': 480}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100000; Y = 8'b11110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2926,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110101; Y = 8'b10011010; // Expected: {'Z': -5406}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110101; Y = 8'b10011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2927,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5406
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001111; Y = 8'b01110100; // Expected: {'Z': -13108}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001111; Y = 8'b01110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2928,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -13108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110001; Y = 8'b11111111; // Expected: {'Z': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110001; Y = 8'b11111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2929,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111001; Y = 8'b00100111; // Expected: {'Z': 4719}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111001; Y = 8'b00100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2930,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4719
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011000; Y = 8'b10010111; // Expected: {'Z': 10920}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011000; Y = 8'b10010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2931,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000111; Y = 8'b01001111; // Expected: {'Z': -9559}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000111; Y = 8'b01001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2932,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9559
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011011; Y = 8'b00001111; // Expected: {'Z': 405}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011011; Y = 8'b00001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2933,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 405
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b00001111; // Expected: {'Z': 915}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b00001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2934,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 915
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100011; Y = 8'b11010000; // Expected: {'Z': -4752}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100011; Y = 8'b11010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2935,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4752
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111100; Y = 8'b00100111; // Expected: {'Z': 4836}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111100; Y = 8'b00100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2936,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4836
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010101; Y = 8'b01001001; // Expected: {'Z': -7811}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010101; Y = 8'b01001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2937,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7811
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010111; Y = 8'b00111010; // Expected: {'Z': 5046}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010111; Y = 8'b00111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2938,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5046
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100000; Y = 8'b11001111; // Expected: {'Z': 4704}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100000; Y = 8'b11001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2939,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4704
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010001; Y = 8'b10111111; // Expected: {'Z': -5265}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010001; Y = 8'b10111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2940,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5265
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b10101110; // Expected: {'Z': -5904}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b10101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2941,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5904
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010111; Y = 8'b00011101; // Expected: {'Z': -1189}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010111; Y = 8'b00011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2942,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110101; Y = 8'b01010100; // Expected: {'Z': 9828}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110101; Y = 8'b01010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2943,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b10111000; // Expected: {'Z': -4896}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b10111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2944,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000001; Y = 8'b10000011; // Expected: {'Z': 15875}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000001; Y = 8'b10000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2945,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 15875
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000100; Y = 8'b10111010; // Expected: {'Z': 4200}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000100; Y = 8'b10111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2946,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111111; Y = 8'b01110111; // Expected: {'Z': -7735}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111111; Y = 8'b01110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2947,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7735
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111100; Y = 8'b00111111; // Expected: {'Z': 3780}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111100; Y = 8'b00111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2948,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111111; Y = 8'b00110011; // Expected: {'Z': -51}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111111; Y = 8'b00110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2949,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011011; Y = 8'b01111010; // Expected: {'Z': -12322}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011011; Y = 8'b01111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2950,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -12322
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010011; Y = 8'b10101011; // Expected: {'Z': 3825}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010011; Y = 8'b10101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2951,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3825
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b11100101; // Expected: {'Z': 2268}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b11100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2952,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2268
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111100; Y = 8'b10010101; // Expected: {'Z': -6420}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111100; Y = 8'b10010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2953,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111110; Y = 8'b11000101; // Expected: {'Z': 118}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111110; Y = 8'b11000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2954,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000111; Y = 8'b11000110; // Expected: {'Z': 3306}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000111; Y = 8'b11000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2955,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3306
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010101; Y = 8'b01111001; // Expected: {'Z': -5203}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010101; Y = 8'b01111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2956,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5203
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111111; Y = 8'b01000001; // Expected: {'Z': 8255}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111111; Y = 8'b01000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2957,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011010; Y = 8'b11010101; // Expected: {'Z': -3870}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011010; Y = 8'b11010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2958,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3870
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010100; Y = 8'b01100111; // Expected: {'Z': 2060}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010100; Y = 8'b01100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2959,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011001; Y = 8'b01100101; // Expected: {'Z': 2525}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011001; Y = 8'b01100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2960,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2525
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111111; Y = 8'b01101111; // Expected: {'Z': 6993}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111111; Y = 8'b01101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2961,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6993
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111101; Y = 8'b01011011; // Expected: {'Z': 11375}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111101; Y = 8'b01011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2962,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11375
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100010; Y = 8'b01100100; // Expected: {'Z': 9800}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100010; Y = 8'b01100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2963,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b11100100; // Expected: {'Z': -532}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b11100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2964,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -532
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b10101000; // Expected: {'Z': -9064}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b10101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2965,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9064
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010111; Y = 8'b00010010; // Expected: {'Z': 1566}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010111; Y = 8'b00010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2966,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1566
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b11110001; // Expected: {'Z': -1845}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b11110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2967,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1845
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100011; Y = 8'b11010101; // Expected: {'Z': -4257}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100011; Y = 8'b11010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2968,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4257
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010101; Y = 8'b00100011; // Expected: {'Z': -1505}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010101; Y = 8'b00100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2969,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1505
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101111; Y = 8'b10110011; // Expected: {'Z': -8547}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101111; Y = 8'b10110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2970,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8547
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b01101110; // Expected: {'Z': -5610}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b01101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2971,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5610
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b00011111; // Expected: {'Z': -1581}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b00011111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2972,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1581
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110111; Y = 8'b10101111; // Expected: {'Z': -9639}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110111; Y = 8'b10101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2973,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9639
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110101; Y = 8'b10001101; // Expected: {'Z': 1265}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110101; Y = 8'b10001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2974,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1265
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111111; Y = 8'b10111110; // Expected: {'Z': 66}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111111; Y = 8'b10111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2975,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100010; Y = 8'b00101111; // Expected: {'Z': -4418}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100010; Y = 8'b00101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2976,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4418
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101000; Y = 8'b01000011; // Expected: {'Z': -5896}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101000; Y = 8'b01000011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2977,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000100; Y = 8'b01101101; // Expected: {'Z': -6540}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000100; Y = 8'b01101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2978,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010010; Y = 8'b10111100; // Expected: {'Z': -1224}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010010; Y = 8'b10111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2979,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111000; Y = 8'b01000101; // Expected: {'Z': 8280}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111000; Y = 8'b01000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2980,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011010; Y = 8'b00001000; // Expected: {'Z': -304}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011010; Y = 8'b00001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2981,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -304
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111000; Y = 8'b01000000; // Expected: {'Z': 3584}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111000; Y = 8'b01000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2982,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3584
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100001; Y = 8'b00010001; // Expected: {'Z': -1615}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100001; Y = 8'b00010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2983,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1615
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b10001000; // Expected: {'Z': -5280}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b10001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2984,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101100; Y = 8'b11101111; // Expected: {'Z': -1836}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101100; Y = 8'b11101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2985,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1836
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001110; Y = 8'b11110100; // Expected: {'Z': -168}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001110; Y = 8'b11110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2986,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100110; Y = 8'b01111010; // Expected: {'Z': 4636}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100110; Y = 8'b01111010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2987,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4636
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010011; Y = 8'b00111111; // Expected: {'Z': 5229}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010011; Y = 8'b00111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2988,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5229
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011000; Y = 8'b10000010; // Expected: {'Z': 13104}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011000; Y = 8'b10000010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2989,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 13104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011001; Y = 8'b11010110; // Expected: {'Z': 4326}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011001; Y = 8'b11010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2990,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4326
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000011; Y = 8'b01010010; // Expected: {'Z': 246}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000011; Y = 8'b01010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2991,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010001; Y = 8'b00111110; // Expected: {'Z': -2914}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010001; Y = 8'b00111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2992,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2914
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b10001110; // Expected: {'Z': 9348}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b10001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2993,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9348
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110110; Y = 8'b01111100; // Expected: {'Z': -1240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110110; Y = 8'b01111100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2994,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111001; Y = 8'b10110000; // Expected: {'Z': -9680}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111001; Y = 8'b10110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2995,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101001; Y = 8'b00001011; // Expected: {'Z': 451}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101001; Y = 8'b00001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2996,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 451
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b01101001; // Expected: {'Z': 4620}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b01101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2997,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111111; Y = 8'b00101010; // Expected: {'Z': 2646}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111111; Y = 8'b00101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2998,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2646
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b00110001; // Expected: {'Z': 98}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b00110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 2999,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011001; Y = 8'b11001100; // Expected: {'Z': -1300}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011001; Y = 8'b11001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3000,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010100; Y = 8'b10001010; // Expected: {'Z': -2360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010100; Y = 8'b10001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3001,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001111; Y = 8'b00100100; // Expected: {'Z': -4068}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001111; Y = 8'b00100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3002,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4068
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010101; Y = 8'b01111111; // Expected: {'Z': 10795}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010101; Y = 8'b01111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3003,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10795
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011000; Y = 8'b00100011; // Expected: {'Z': 840}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011000; Y = 8'b00100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3004,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b10111101; // Expected: {'Z': -7504}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b10111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3005,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000011; Y = 8'b10110000; // Expected: {'Z': -240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000011; Y = 8'b10110000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3006,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011111; Y = 8'b00001001; // Expected: {'Z': -297}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011111; Y = 8'b00001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3007,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -297
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110010; Y = 8'b10000100; // Expected: {'Z': -6200}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110010; Y = 8'b10000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3008,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b01111101; // Expected: {'Z': 750}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b01111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3009,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101001; Y = 8'b01100111; // Expected: {'Z': -2369}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101001; Y = 8'b01100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3010,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2369
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100101; Y = 8'b10101101; // Expected: {'Z': 2241}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100101; Y = 8'b10101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3011,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010001; Y = 8'b11101110; // Expected: {'Z': 846}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010001; Y = 8'b11101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3012,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 846
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b00001111; // Expected: {'Z': 225}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b00001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3013,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110010; Y = 8'b01010101; // Expected: {'Z': -6630}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110010; Y = 8'b01010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3014,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6630
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111011; Y = 8'b00100000; // Expected: {'Z': -2208}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111011; Y = 8'b00100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3015,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001111; Y = 8'b01101110; // Expected: {'Z': -5390}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001111; Y = 8'b01101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3016,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5390
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001000; Y = 8'b10111011; // Expected: {'Z': -552}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001000; Y = 8'b10111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3017,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001111; Y = 8'b11011110; // Expected: {'Z': 1666}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001111; Y = 8'b11011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3018,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1666
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011001; Y = 8'b01111011; // Expected: {'Z': 10947}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011001; Y = 8'b01111011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3019,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 10947
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010100; Y = 8'b10010110; // Expected: {'Z': -2120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010100; Y = 8'b10010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3020,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101011; Y = 8'b01010111; // Expected: {'Z': 9309}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101011; Y = 8'b01010111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3021,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9309
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101100; Y = 8'b01111110; // Expected: {'Z': 13608}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101100; Y = 8'b01111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3022,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 13608
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101100; Y = 8'b11001001; // Expected: {'Z': -5940}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101100; Y = 8'b11001001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3023,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5940
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000011; Y = 8'b00010000; // Expected: {'Z': 48}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000011; Y = 8'b00010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3024,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101011; Y = 8'b10110100; // Expected: {'Z': -3268}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00101011; Y = 8'b10110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3025,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3268
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010110; Y = 8'b11011000; // Expected: {'Z': -3440}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010110; Y = 8'b11011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3026,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111000; Y = 8'b00101100; // Expected: {'Z': -352}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111000; Y = 8'b00101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3027,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001001; Y = 8'b00011000; // Expected: {'Z': -1320}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001001; Y = 8'b00011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3028,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001110; Y = 8'b11001010; // Expected: {'Z': 6156}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001110; Y = 8'b11001010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3029,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010000; Y = 8'b11010000; // Expected: {'Z': -3840}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010000; Y = 8'b11010000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3030,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110001; Y = 8'b01001101; // Expected: {'Z': -1155}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110001; Y = 8'b01001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3031,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b11000000; // Expected: {'Z': -384}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b11000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3032,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -384
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100000; Y = 8'b10111111; // Expected: {'Z': 6240}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100000; Y = 8'b10111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3033,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111000; Y = 8'b11110111; // Expected: {'Z': -504}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111000; Y = 8'b11110111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3034,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111101; Y = 8'b10010101; // Expected: {'Z': 321}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111101; Y = 8'b10010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3035,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 321
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101101; Y = 8'b11010001; // Expected: {'Z': 893}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101101; Y = 8'b11010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3036,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 893
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011011; Y = 8'b11101011; // Expected: {'Z': -567}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011011; Y = 8'b11101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3037,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -567
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b00100111; // Expected: {'Z': 858}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b00100111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3038,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 858
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000110; Y = 8'b11111111; // Expected: {'Z': -70}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000110; Y = 8'b11111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3039,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110011; Y = 8'b11100000; // Expected: {'Z': -1632}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110011; Y = 8'b11100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3040,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1632
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110001; Y = 8'b00100011; // Expected: {'Z': -525}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110001; Y = 8'b00100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3041,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -525
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100100; Y = 8'b11110110; // Expected: {'Z': 920}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100100; Y = 8'b11110110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3042,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b00100100; // Expected: {'Z': 3168}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b00100100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3043,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011010; Y = 8'b10100001; // Expected: {'Z': -8550}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011010; Y = 8'b10100001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3044,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100101; Y = 8'b00001000; // Expected: {'Z': -216}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11100101; Y = 8'b00001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3045,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b01010011; // Expected: {'Z': 4482}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b01010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3046,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4482
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111000; Y = 8'b00011100; // Expected: {'Z': 1568}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111000; Y = 8'b00011100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3047,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1568
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b11000001; // Expected: {'Z': -4284}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b11000001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3048,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4284
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b10110010; // Expected: {'Z': 4368}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b10110010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3049,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011011; Y = 8'b01111111; // Expected: {'Z': -4699}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011011; Y = 8'b01111111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3050,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4699
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000100; Y = 8'b10101111; // Expected: {'Z': 4860}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000100; Y = 8'b10101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3051,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4860
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100001; Y = 8'b01101100; // Expected: {'Z': -10260}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100001; Y = 8'b01101100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3052,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -10260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b10101110; // Expected: {'Z': -5904}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b10101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3053,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -5904
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001100; Y = 8'b01010110; // Expected: {'Z': -9976}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10001100; Y = 8'b01010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3054,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9976
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011100; Y = 8'b00010110; // Expected: {'Z': 2024}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011100; Y = 8'b00010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3055,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011110; Y = 8'b01001011; // Expected: {'Z': -2550}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011110; Y = 8'b01001011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3056,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b11100110; // Expected: {'Z': -2496}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b11100110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3057,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100011; Y = 8'b10101101; // Expected: {'Z': 7719}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10100011; Y = 8'b10101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3058,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7719
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b11011001; // Expected: {'Z': -3744}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b11011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3059,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3744
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001110; Y = 8'b01111110; // Expected: {'Z': 1764}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001110; Y = 8'b01111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3060,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1764
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b01101000; // Expected: {'Z': -6136}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b01101000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3061,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010011; Y = 8'b10010011; // Expected: {'Z': -9047}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01010011; Y = 8'b10010011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3062,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9047
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010111; Y = 8'b10110100; // Expected: {'Z': 7980}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010111; Y = 8'b10110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3063,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 7980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000100; Y = 8'b00011101; // Expected: {'Z': -1740}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000100; Y = 8'b00011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3064,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1740
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111001; Y = 8'b11110100; // Expected: {'Z': 84}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11111001; Y = 8'b11110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3065,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011100; Y = 8'b11111001; // Expected: {'Z': -196}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011100; Y = 8'b11111001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3066,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b10101111; // Expected: {'Z': -8343}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b10101111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3067,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8343
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101100; Y = 8'b01000110; // Expected: {'Z': -1400}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101100; Y = 8'b01000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3068,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110101; Y = 8'b11100000; // Expected: {'Z': 352}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110101; Y = 8'b11100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3069,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111011; Y = 8'b01110001; // Expected: {'Z': -7797}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111011; Y = 8'b01110001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3070,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -7797
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000000; Y = 8'b11000101; // Expected: {'Z': -3776}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01000000; Y = 8'b11000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3071,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3776
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101101; Y = 8'b00000100; // Expected: {'Z': 436}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01101101; Y = 8'b00000100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3072,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 436
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010111; Y = 8'b00100000; // Expected: {'Z': -3360}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010111; Y = 8'b00100000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3073,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001010; Y = 8'b11001100; // Expected: {'Z': 2808}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001010; Y = 8'b11001100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3074,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011010; Y = 8'b01011001; // Expected: {'Z': 8010}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011010; Y = 8'b01011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3075,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8010
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b01111000; // Expected: {'Z': -6120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b01111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3076,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b10001111; // Expected: {'Z': -1695}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b10001111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3077,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1695
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001001; Y = 8'b00000111; // Expected: {'Z': -385}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11001001; Y = 8'b00000111; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3078,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -385
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011101; Y = 8'b00101001; // Expected: {'Z': -4059}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011101; Y = 8'b00101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3079,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -4059
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000000; Y = 8'b10101001; // Expected: {'Z': 11136}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10000000; Y = 8'b10101001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3080,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 11136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011101; Y = 8'b01011011; // Expected: {'Z': 8463}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011101; Y = 8'b01011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3081,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 8463
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110001; Y = 8'b01010101; // Expected: {'Z': 9605}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01110001; Y = 8'b01010101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3082,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 9605
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110111; Y = 8'b01001000; // Expected: {'Z': -648}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11110111; Y = 8'b01001000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3083,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100001; Y = 8'b00101110; // Expected: {'Z': 4462}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100001; Y = 8'b00101110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3084,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b00001110; // Expected: {'Z': 84}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b00001110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3085,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b01011011; // Expected: {'Z': 819}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b01011011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3086,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 819
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101101; Y = 8'b11100011; // Expected: {'Z': 551}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101101; Y = 8'b11100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3087,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 551
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111000; Y = 8'b01011001; // Expected: {'Z': -6408}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111000; Y = 8'b01011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3088,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b10111000; // Expected: {'Z': 4248}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b10111000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3089,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110010; Y = 8'b00000110; // Expected: {'Z': -468}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110010; Y = 8'b00000110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3090,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -468
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b01000000; // Expected: {'Z': 6144}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b01000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3091,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b10111110; // Expected: {'Z': -2376}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b10111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3092,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -2376
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111110; Y = 8'b10110011; // Expected: {'Z': -9702}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01111110; Y = 8'b10110011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3093,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -9702
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101011; Y = 8'b11011110; // Expected: {'Z': 714}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11101011; Y = 8'b11011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3094,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 714
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110111; Y = 8'b11011101; // Expected: {'Z': -1925}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00110111; Y = 8'b11011101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3095,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1925
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011011; Y = 8'b11101101; // Expected: {'Z': -513}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011011; Y = 8'b11101101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3096,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -513
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101010; Y = 8'b10110101; // Expected: {'Z': 6450}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101010; Y = 8'b10110101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3097,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 6450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011011; Y = 8'b10000101; // Expected: {'Z': 4551}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011011; Y = 8'b10000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3098,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4551
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000000; Y = 8'b00111101; // Expected: {'Z': -3904}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11000000; Y = 8'b00111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3099,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3904
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011101; Y = 8'b00101010; // Expected: {'Z': -1470}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11011101; Y = 8'b00101010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3100,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1470
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110100; Y = 8'b00101011; // Expected: {'Z': -3268}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110100; Y = 8'b00101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3101,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -3268
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011111; Y = 8'b01100011; // Expected: {'Z': 3069}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011111; Y = 8'b01100011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3102,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 3069
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101111; Y = 8'b01010001; // Expected: {'Z': -6561}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10101111; Y = 8'b01010001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3103,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -6561
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100010; Y = 8'b00101011; // Expected: {'Z': 4214}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01100010; Y = 8'b00101011; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3104,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111111; Y = 8'b01010110; // Expected: {'Z': 5418}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00111111; Y = 8'b01010110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3105,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5418
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011011; Y = 8'b00011010; // Expected: {'Z': 2366}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011011; Y = 8'b00011010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3106,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2366
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b11010100; // Expected: {'Z': -572}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b11010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3107,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -572
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000100; Y = 8'b11100101; // Expected: {'Z': -108}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00000100; Y = 8'b11100101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3108,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110111; Y = 8'b11111101; // Expected: {'Z': 219}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110111; Y = 8'b11111101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3109,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 219
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010010; Y = 8'b00011000; // Expected: {'Z': 432}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00010010; Y = 8'b00011000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3110,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b00000000; // Expected: {'Z': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b00000000; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3111,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011101; Y = 8'b01011001; // Expected: {'Z': -8811}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011101; Y = 8'b01011001; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3112,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -8811
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110000; Y = 8'b00000101; // Expected: {'Z': -400}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10110000; Y = 8'b00000101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3113,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010011; Y = 8'b11010100; // Expected: {'Z': 4796}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010011; Y = 8'b11010100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3114,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4796
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111000; Y = 8'b00010010; // Expected: {'Z': -1296}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111000; Y = 8'b00010010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3115,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111001; Y = 8'b11100010; // Expected: {'Z': 2130}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10111001; Y = 8'b11100010; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3116,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 2130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010011; Y = 8'b10011110; // Expected: {'Z': 4410}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b11010011; Y = 8'b10011110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3117,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4410
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001100; Y = 8'b00111110; // Expected: {'Z': 4712}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b01001100; Y = 8'b00111110; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3118,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 4712
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b11001101; // Expected: {'Z': -1479}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b11001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3119,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 -1479
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010010; Y = 8'b11110100; // Expected: {'Z': 1320}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10010010; Y = 8'b11110100; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3120,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 1320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011000; Y = 8'b11001101; // Expected: {'Z': 5304}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        wait(~valid);
        
        $display("Test %0d: Inputs: X = 8'b10011000; Y = 8'b11001101; | Outputs: Z=%b, valid=%b | Expected: Z=%d",
                 3121,
                 
                 Z, 
                 
                 valid
                 , 
                 
                 5304
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        $finish;
    end
  
endmodule