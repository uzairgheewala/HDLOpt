
`timescale 1ns / 1ps

module tb_N8_array_multiplier;

    // Parameters
    
    parameter N = 8;
    
     
    // Inputs
    
    reg  [7:0] A;
    
    reg  [7:0] B;
    
    
    // Outputs
    
    wire   P;
    
    
    // Instantiate the Unit Under Test (UUT)
    array_multiplier  #( N ) uut (
        
        .A(A),
        
        .B(B),
        
        
        .P(P)
        
    );

    // Clock generation 
    

    
    
    initial begin
        // Initialize Inputs
        
        A = 0;
        
        B = 0;
        
    
        // Wait for global reset
        #100;
    
        // Stimuli
        
        #10 A = 8'b10001110; B = 8'b11000101; // Expected: {'P': 27974}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001110; B = 8'b11000101; | Outputs: P=%b | Expected: P=%d",
                 0,
                 
                 P
                 , 
                 
                 27974
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001000; B = 8'b01111001; // Expected: {'P': 968}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001000; B = 8'b01111001; | Outputs: P=%b | Expected: P=%d",
                 1,
                 
                 P
                 , 
                 
                 968
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000011; B = 8'b01011110; // Expected: {'P': 282}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000011; B = 8'b01011110; | Outputs: P=%b | Expected: P=%d",
                 2,
                 
                 P
                 , 
                 
                 282
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110010; B = 8'b01010101; // Expected: {'P': 20570}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110010; B = 8'b01010101; | Outputs: P=%b | Expected: P=%d",
                 3,
                 
                 P
                 , 
                 
                 20570
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100010; B = 8'b01000010; // Expected: {'P': 6468}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100010; B = 8'b01000010; | Outputs: P=%b | Expected: P=%d",
                 4,
                 
                 P
                 , 
                 
                 6468
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101010; B = 8'b00010110; // Expected: {'P': 5148}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101010; B = 8'b00010110; | Outputs: P=%b | Expected: P=%d",
                 5,
                 
                 P
                 , 
                 
                 5148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101010; B = 8'b11011111; // Expected: {'P': 23638}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101010; B = 8'b11011111; | Outputs: P=%b | Expected: P=%d",
                 6,
                 
                 P
                 , 
                 
                 23638
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011110; B = 8'b11101110; // Expected: {'P': 22372}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011110; B = 8'b11101110; | Outputs: P=%b | Expected: P=%d",
                 7,
                 
                 P
                 , 
                 
                 22372
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110101; B = 8'b11011011; // Expected: {'P': 25623}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110101; B = 8'b11011011; | Outputs: P=%b | Expected: P=%d",
                 8,
                 
                 P
                 , 
                 
                 25623
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000010; B = 8'b01110110; // Expected: {'P': 22892}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000010; B = 8'b01110110; | Outputs: P=%b | Expected: P=%d",
                 9,
                 
                 P
                 , 
                 
                 22892
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000100; B = 8'b10111110; // Expected: {'P': 25080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000100; B = 8'b10111110; | Outputs: P=%b | Expected: P=%d",
                 10,
                 
                 P
                 , 
                 
                 25080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110100; B = 8'b11011000; // Expected: {'P': 11232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110100; B = 8'b11011000; | Outputs: P=%b | Expected: P=%d",
                 11,
                 
                 P
                 , 
                 
                 11232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110010; B = 8'b01010101; // Expected: {'P': 9690}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110010; B = 8'b01010101; | Outputs: P=%b | Expected: P=%d",
                 12,
                 
                 P
                 , 
                 
                 9690
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010101; B = 8'b01110011; // Expected: {'P': 24495}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010101; B = 8'b01110011; | Outputs: P=%b | Expected: P=%d",
                 13,
                 
                 P
                 , 
                 
                 24495
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011100; B = 8'b11001010; // Expected: {'P': 31512}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011100; B = 8'b11001010; | Outputs: P=%b | Expected: P=%d",
                 14,
                 
                 P
                 , 
                 
                 31512
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001101; B = 8'b01010001; // Expected: {'P': 6237}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001101; B = 8'b01010001; | Outputs: P=%b | Expected: P=%d",
                 15,
                 
                 P
                 , 
                 
                 6237
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000011; B = 8'b00110100; // Expected: {'P': 3484}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000011; B = 8'b00110100; | Outputs: P=%b | Expected: P=%d",
                 16,
                 
                 P
                 , 
                 
                 3484
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000011; B = 8'b11111100; // Expected: {'P': 49140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000011; B = 8'b11111100; | Outputs: P=%b | Expected: P=%d",
                 17,
                 
                 P
                 , 
                 
                 49140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000100; B = 8'b10000111; // Expected: {'P': 17820}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000100; B = 8'b10000111; | Outputs: P=%b | Expected: P=%d",
                 18,
                 
                 P
                 , 
                 
                 17820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111010; B = 8'b10001000; // Expected: {'P': 34000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111010; B = 8'b10001000; | Outputs: P=%b | Expected: P=%d",
                 19,
                 
                 P
                 , 
                 
                 34000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001101; B = 8'b10011001; // Expected: {'P': 1989}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001101; B = 8'b10011001; | Outputs: P=%b | Expected: P=%d",
                 20,
                 
                 P
                 , 
                 
                 1989
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010001; B = 8'b11010010; // Expected: {'P': 30450}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010001; B = 8'b11010010; | Outputs: P=%b | Expected: P=%d",
                 21,
                 
                 P
                 , 
                 
                 30450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111100; B = 8'b10101101; // Expected: {'P': 32524}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111100; B = 8'b10101101; | Outputs: P=%b | Expected: P=%d",
                 22,
                 
                 P
                 , 
                 
                 32524
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111100; B = 8'b10000110; // Expected: {'P': 33768}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111100; B = 8'b10000110; | Outputs: P=%b | Expected: P=%d",
                 23,
                 
                 P
                 , 
                 
                 33768
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101100; B = 8'b01110111; // Expected: {'P': 20468}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101100; B = 8'b01110111; | Outputs: P=%b | Expected: P=%d",
                 24,
                 
                 P
                 , 
                 
                 20468
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010111; B = 8'b10111001; // Expected: {'P': 27935}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010111; B = 8'b10111001; | Outputs: P=%b | Expected: P=%d",
                 25,
                 
                 P
                 , 
                 
                 27935
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101001; B = 8'b11010000; // Expected: {'P': 8528}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101001; B = 8'b11010000; | Outputs: P=%b | Expected: P=%d",
                 26,
                 
                 P
                 , 
                 
                 8528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000100; B = 8'b11011101; // Expected: {'P': 43316}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000100; B = 8'b11011101; | Outputs: P=%b | Expected: P=%d",
                 27,
                 
                 P
                 , 
                 
                 43316
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110100; B = 8'b00010001; // Expected: {'P': 4148}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110100; B = 8'b00010001; | Outputs: P=%b | Expected: P=%d",
                 28,
                 
                 P
                 , 
                 
                 4148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110100; B = 8'b11000111; // Expected: {'P': 10348}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110100; B = 8'b11000111; | Outputs: P=%b | Expected: P=%d",
                 29,
                 
                 P
                 , 
                 
                 10348
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111100; B = 8'b01001101; // Expected: {'P': 19404}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111100; B = 8'b01001101; | Outputs: P=%b | Expected: P=%d",
                 30,
                 
                 P
                 , 
                 
                 19404
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100111; B = 8'b10010011; // Expected: {'P': 24549}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100111; B = 8'b10010011; | Outputs: P=%b | Expected: P=%d",
                 31,
                 
                 P
                 , 
                 
                 24549
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011100; B = 8'b10010010; // Expected: {'P': 32120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011100; B = 8'b10010010; | Outputs: P=%b | Expected: P=%d",
                 32,
                 
                 P
                 , 
                 
                 32120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000000; B = 8'b10110110; // Expected: {'P': 23296}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000000; B = 8'b10110110; | Outputs: P=%b | Expected: P=%d",
                 33,
                 
                 P
                 , 
                 
                 23296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110011; B = 8'b01001000; // Expected: {'P': 17496}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110011; B = 8'b01001000; | Outputs: P=%b | Expected: P=%d",
                 34,
                 
                 P
                 , 
                 
                 17496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001110; B = 8'b00111110; // Expected: {'P': 8804}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001110; B = 8'b00111110; | Outputs: P=%b | Expected: P=%d",
                 35,
                 
                 P
                 , 
                 
                 8804
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011111; B = 8'b10010001; // Expected: {'P': 23055}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011111; B = 8'b10010001; | Outputs: P=%b | Expected: P=%d",
                 36,
                 
                 P
                 , 
                 
                 23055
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001100; B = 8'b01011010; // Expected: {'P': 18360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001100; B = 8'b01011010; | Outputs: P=%b | Expected: P=%d",
                 37,
                 
                 P
                 , 
                 
                 18360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010110; B = 8'b11011001; // Expected: {'P': 46438}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010110; B = 8'b11011001; | Outputs: P=%b | Expected: P=%d",
                 38,
                 
                 P
                 , 
                 
                 46438
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110111; B = 8'b01010100; // Expected: {'P': 9996}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110111; B = 8'b01010100; | Outputs: P=%b | Expected: P=%d",
                 39,
                 
                 P
                 , 
                 
                 9996
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010010; B = 8'b01111001; // Expected: {'P': 17666}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010010; B = 8'b01111001; | Outputs: P=%b | Expected: P=%d",
                 40,
                 
                 P
                 , 
                 
                 17666
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100011; B = 8'b10110100; // Expected: {'P': 40860}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100011; B = 8'b10110100; | Outputs: P=%b | Expected: P=%d",
                 41,
                 
                 P
                 , 
                 
                 40860
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011110; B = 8'b10010110; // Expected: {'P': 33300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011110; B = 8'b10010110; | Outputs: P=%b | Expected: P=%d",
                 42,
                 
                 P
                 , 
                 
                 33300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011001; B = 8'b10010010; // Expected: {'P': 12994}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011001; B = 8'b10010010; | Outputs: P=%b | Expected: P=%d",
                 43,
                 
                 P
                 , 
                 
                 12994
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101000; B = 8'b00001001; // Expected: {'P': 1512}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101000; B = 8'b00001001; | Outputs: P=%b | Expected: P=%d",
                 44,
                 
                 P
                 , 
                 
                 1512
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000110; B = 8'b11101010; // Expected: {'P': 46332}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000110; B = 8'b11101010; | Outputs: P=%b | Expected: P=%d",
                 45,
                 
                 P
                 , 
                 
                 46332
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001011; B = 8'b11001000; // Expected: {'P': 15000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001011; B = 8'b11001000; | Outputs: P=%b | Expected: P=%d",
                 46,
                 
                 P
                 , 
                 
                 15000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011100; B = 8'b01010000; // Expected: {'P': 7360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011100; B = 8'b01010000; | Outputs: P=%b | Expected: P=%d",
                 47,
                 
                 P
                 , 
                 
                 7360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101000; B = 8'b11010000; // Expected: {'P': 48256}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101000; B = 8'b11010000; | Outputs: P=%b | Expected: P=%d",
                 48,
                 
                 P
                 , 
                 
                 48256
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100101; B = 8'b11110100; // Expected: {'P': 40260}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100101; B = 8'b11110100; | Outputs: P=%b | Expected: P=%d",
                 49,
                 
                 P
                 , 
                 
                 40260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010100; B = 8'b00001010; // Expected: {'P': 840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010100; B = 8'b00001010; | Outputs: P=%b | Expected: P=%d",
                 50,
                 
                 P
                 , 
                 
                 840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011011; B = 8'b01000111; // Expected: {'P': 1917}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011011; B = 8'b01000111; | Outputs: P=%b | Expected: P=%d",
                 51,
                 
                 P
                 , 
                 
                 1917
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010010; B = 8'b11110011; // Expected: {'P': 51030}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010010; B = 8'b11110011; | Outputs: P=%b | Expected: P=%d",
                 52,
                 
                 P
                 , 
                 
                 51030
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111000; B = 8'b11010111; // Expected: {'P': 53320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111000; B = 8'b11010111; | Outputs: P=%b | Expected: P=%d",
                 53,
                 
                 P
                 , 
                 
                 53320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011101; B = 8'b01110100; // Expected: {'P': 18212}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011101; B = 8'b01110100; | Outputs: P=%b | Expected: P=%d",
                 54,
                 
                 P
                 , 
                 
                 18212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100110; B = 8'b01000110; // Expected: {'P': 2660}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100110; B = 8'b01000110; | Outputs: P=%b | Expected: P=%d",
                 55,
                 
                 P
                 , 
                 
                 2660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100111; B = 8'b10011010; // Expected: {'P': 6006}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100111; B = 8'b10011010; | Outputs: P=%b | Expected: P=%d",
                 56,
                 
                 P
                 , 
                 
                 6006
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100010; B = 8'b00111101; // Expected: {'P': 13786}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100010; B = 8'b00111101; | Outputs: P=%b | Expected: P=%d",
                 57,
                 
                 P
                 , 
                 
                 13786
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110100; B = 8'b00010100; // Expected: {'P': 4880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110100; B = 8'b00010100; | Outputs: P=%b | Expected: P=%d",
                 58,
                 
                 P
                 , 
                 
                 4880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110000; B = 8'b11101101; // Expected: {'P': 26544}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110000; B = 8'b11101101; | Outputs: P=%b | Expected: P=%d",
                 59,
                 
                 P
                 , 
                 
                 26544
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110111; B = 8'b10001100; // Expected: {'P': 16660}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110111; B = 8'b10001100; | Outputs: P=%b | Expected: P=%d",
                 60,
                 
                 P
                 , 
                 
                 16660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111110; B = 8'b11001111; // Expected: {'P': 26082}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111110; B = 8'b11001111; | Outputs: P=%b | Expected: P=%d",
                 61,
                 
                 P
                 , 
                 
                 26082
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100011; B = 8'b01001011; // Expected: {'P': 7425}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100011; B = 8'b01001011; | Outputs: P=%b | Expected: P=%d",
                 62,
                 
                 P
                 , 
                 
                 7425
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110010; B = 8'b11111110; // Expected: {'P': 28956}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110010; B = 8'b11111110; | Outputs: P=%b | Expected: P=%d",
                 63,
                 
                 P
                 , 
                 
                 28956
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101001; B = 8'b01101110; // Expected: {'P': 25630}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101001; B = 8'b01101110; | Outputs: P=%b | Expected: P=%d",
                 64,
                 
                 P
                 , 
                 
                 25630
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110011; B = 8'b01010001; // Expected: {'P': 4131}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110011; B = 8'b01010001; | Outputs: P=%b | Expected: P=%d",
                 65,
                 
                 P
                 , 
                 
                 4131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010110; B = 8'b10110000; // Expected: {'P': 3872}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010110; B = 8'b10110000; | Outputs: P=%b | Expected: P=%d",
                 66,
                 
                 P
                 , 
                 
                 3872
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101110; B = 8'b00111010; // Expected: {'P': 13804}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101110; B = 8'b00111010; | Outputs: P=%b | Expected: P=%d",
                 67,
                 
                 P
                 , 
                 
                 13804
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001001; B = 8'b00011111; // Expected: {'P': 2263}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001001; B = 8'b00011111; | Outputs: P=%b | Expected: P=%d",
                 68,
                 
                 P
                 , 
                 
                 2263
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001010; B = 8'b10111010; // Expected: {'P': 1860}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001010; B = 8'b10111010; | Outputs: P=%b | Expected: P=%d",
                 69,
                 
                 P
                 , 
                 
                 1860
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010011; B = 8'b11010000; // Expected: {'P': 30576}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010011; B = 8'b11010000; | Outputs: P=%b | Expected: P=%d",
                 70,
                 
                 P
                 , 
                 
                 30576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011101; B = 8'b01001111; // Expected: {'P': 17459}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011101; B = 8'b01001111; | Outputs: P=%b | Expected: P=%d",
                 71,
                 
                 P
                 , 
                 
                 17459
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111000; B = 8'b10011001; // Expected: {'P': 18360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111000; B = 8'b10011001; | Outputs: P=%b | Expected: P=%d",
                 72,
                 
                 P
                 , 
                 
                 18360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111101; B = 8'b01110100; // Expected: {'P': 14500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111101; B = 8'b01110100; | Outputs: P=%b | Expected: P=%d",
                 73,
                 
                 P
                 , 
                 
                 14500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001011; B = 8'b00001101; // Expected: {'P': 975}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001011; B = 8'b00001101; | Outputs: P=%b | Expected: P=%d",
                 74,
                 
                 P
                 , 
                 
                 975
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100101; B = 8'b10110010; // Expected: {'P': 6586}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100101; B = 8'b10110010; | Outputs: P=%b | Expected: P=%d",
                 75,
                 
                 P
                 , 
                 
                 6586
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111111; B = 8'b00001011; // Expected: {'P': 2805}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111111; B = 8'b00001011; | Outputs: P=%b | Expected: P=%d",
                 76,
                 
                 P
                 , 
                 
                 2805
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110111; B = 8'b10111101; // Expected: {'P': 46683}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110111; B = 8'b10111101; | Outputs: P=%b | Expected: P=%d",
                 77,
                 
                 P
                 , 
                 
                 46683
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101100; B = 8'b11000111; // Expected: {'P': 46964}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101100; B = 8'b11000111; | Outputs: P=%b | Expected: P=%d",
                 78,
                 
                 P
                 , 
                 
                 46964
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011011; B = 8'b10010110; // Expected: {'P': 4050}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011011; B = 8'b10010110; | Outputs: P=%b | Expected: P=%d",
                 79,
                 
                 P
                 , 
                 
                 4050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101111; B = 8'b01000100; // Expected: {'P': 7548}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101111; B = 8'b01000100; | Outputs: P=%b | Expected: P=%d",
                 80,
                 
                 P
                 , 
                 
                 7548
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111111; B = 8'b01000001; // Expected: {'P': 16575}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111111; B = 8'b01000001; | Outputs: P=%b | Expected: P=%d",
                 81,
                 
                 P
                 , 
                 
                 16575
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011000; B = 8'b10100010; // Expected: {'P': 24624}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011000; B = 8'b10100010; | Outputs: P=%b | Expected: P=%d",
                 82,
                 
                 P
                 , 
                 
                 24624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000100; B = 8'b11110000; // Expected: {'P': 16320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000100; B = 8'b11110000; | Outputs: P=%b | Expected: P=%d",
                 83,
                 
                 P
                 , 
                 
                 16320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001000; B = 8'b00111010; // Expected: {'P': 11600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001000; B = 8'b00111010; | Outputs: P=%b | Expected: P=%d",
                 84,
                 
                 P
                 , 
                 
                 11600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000000; B = 8'b01000000; // Expected: {'P': 12288}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000000; B = 8'b01000000; | Outputs: P=%b | Expected: P=%d",
                 85,
                 
                 P
                 , 
                 
                 12288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000010; B = 8'b00001010; // Expected: {'P': 1300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000010; B = 8'b00001010; | Outputs: P=%b | Expected: P=%d",
                 86,
                 
                 P
                 , 
                 
                 1300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110010; B = 8'b01000011; // Expected: {'P': 11926}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110010; B = 8'b01000011; | Outputs: P=%b | Expected: P=%d",
                 87,
                 
                 P
                 , 
                 
                 11926
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100100; B = 8'b10010101; // Expected: {'P': 5364}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100100; B = 8'b10010101; | Outputs: P=%b | Expected: P=%d",
                 88,
                 
                 P
                 , 
                 
                 5364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111101; B = 8'b00110100; // Expected: {'P': 9828}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111101; B = 8'b00110100; | Outputs: P=%b | Expected: P=%d",
                 89,
                 
                 P
                 , 
                 
                 9828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001001; B = 8'b01001110; // Expected: {'P': 5694}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001001; B = 8'b01001110; | Outputs: P=%b | Expected: P=%d",
                 90,
                 
                 P
                 , 
                 
                 5694
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111010; B = 8'b10101000; // Expected: {'P': 9744}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111010; B = 8'b10101000; | Outputs: P=%b | Expected: P=%d",
                 91,
                 
                 P
                 , 
                 
                 9744
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101111; B = 8'b10110100; // Expected: {'P': 43020}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101111; B = 8'b10110100; | Outputs: P=%b | Expected: P=%d",
                 92,
                 
                 P
                 , 
                 
                 43020
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110001; B = 8'b10001010; // Expected: {'P': 15594}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110001; B = 8'b10001010; | Outputs: P=%b | Expected: P=%d",
                 93,
                 
                 P
                 , 
                 
                 15594
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111100; B = 8'b10101100; // Expected: {'P': 43344}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111100; B = 8'b10101100; | Outputs: P=%b | Expected: P=%d",
                 94,
                 
                 P
                 , 
                 
                 43344
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100101; B = 8'b10100001; // Expected: {'P': 5957}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100101; B = 8'b10100001; | Outputs: P=%b | Expected: P=%d",
                 95,
                 
                 P
                 , 
                 
                 5957
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101010; B = 8'b01100111; // Expected: {'P': 24102}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101010; B = 8'b01100111; | Outputs: P=%b | Expected: P=%d",
                 96,
                 
                 P
                 , 
                 
                 24102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010110; B = 8'b10001011; // Expected: {'P': 20850}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010110; B = 8'b10001011; | Outputs: P=%b | Expected: P=%d",
                 97,
                 
                 P
                 , 
                 
                 20850
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011101; B = 8'b00010111; // Expected: {'P': 3611}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011101; B = 8'b00010111; | Outputs: P=%b | Expected: P=%d",
                 98,
                 
                 P
                 , 
                 
                 3611
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101011; B = 8'b00001000; // Expected: {'P': 856}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101011; B = 8'b00001000; | Outputs: P=%b | Expected: P=%d",
                 99,
                 
                 P
                 , 
                 
                 856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101100; B = 8'b10111000; // Expected: {'P': 31648}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101100; B = 8'b10111000; | Outputs: P=%b | Expected: P=%d",
                 100,
                 
                 P
                 , 
                 
                 31648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101001; B = 8'b10111011; // Expected: {'P': 43571}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101001; B = 8'b10111011; | Outputs: P=%b | Expected: P=%d",
                 101,
                 
                 P
                 , 
                 
                 43571
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111011; B = 8'b10101111; // Expected: {'P': 43925}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111011; B = 8'b10101111; | Outputs: P=%b | Expected: P=%d",
                 102,
                 
                 P
                 , 
                 
                 43925
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100101; B = 8'b10110111; // Expected: {'P': 6771}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100101; B = 8'b10110111; | Outputs: P=%b | Expected: P=%d",
                 103,
                 
                 P
                 , 
                 
                 6771
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101110; B = 8'b01101010; // Expected: {'P': 18444}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101110; B = 8'b01101010; | Outputs: P=%b | Expected: P=%d",
                 104,
                 
                 P
                 , 
                 
                 18444
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100110; B = 8'b10101001; // Expected: {'P': 6422}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100110; B = 8'b10101001; | Outputs: P=%b | Expected: P=%d",
                 105,
                 
                 P
                 , 
                 
                 6422
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001000; B = 8'b00111000; // Expected: {'P': 11200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001000; B = 8'b00111000; | Outputs: P=%b | Expected: P=%d",
                 106,
                 
                 P
                 , 
                 
                 11200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100110; B = 8'b10101011; // Expected: {'P': 17442}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100110; B = 8'b10101011; | Outputs: P=%b | Expected: P=%d",
                 107,
                 
                 P
                 , 
                 
                 17442
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011100; B = 8'b10000010; // Expected: {'P': 3640}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011100; B = 8'b10000010; | Outputs: P=%b | Expected: P=%d",
                 108,
                 
                 P
                 , 
                 
                 3640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001111; B = 8'b01010100; // Expected: {'P': 17388}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001111; B = 8'b01010100; | Outputs: P=%b | Expected: P=%d",
                 109,
                 
                 P
                 , 
                 
                 17388
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101011; B = 8'b01111001; // Expected: {'P': 28435}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101011; B = 8'b01111001; | Outputs: P=%b | Expected: P=%d",
                 110,
                 
                 P
                 , 
                 
                 28435
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001110; B = 8'b01010101; // Expected: {'P': 6630}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001110; B = 8'b01010101; | Outputs: P=%b | Expected: P=%d",
                 111,
                 
                 P
                 , 
                 
                 6630
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011101; B = 8'b10101011; // Expected: {'P': 4959}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011101; B = 8'b10101011; | Outputs: P=%b | Expected: P=%d",
                 112,
                 
                 P
                 , 
                 
                 4959
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100101; B = 8'b00100111; // Expected: {'P': 6435}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100101; B = 8'b00100111; | Outputs: P=%b | Expected: P=%d",
                 113,
                 
                 P
                 , 
                 
                 6435
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010000; B = 8'b01101100; // Expected: {'P': 22464}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010000; B = 8'b01101100; | Outputs: P=%b | Expected: P=%d",
                 114,
                 
                 P
                 , 
                 
                 22464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001010; B = 8'b00000001; // Expected: {'P': 202}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001010; B = 8'b00000001; | Outputs: P=%b | Expected: P=%d",
                 115,
                 
                 P
                 , 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110000; B = 8'b10010100; // Expected: {'P': 35520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110000; B = 8'b10010100; | Outputs: P=%b | Expected: P=%d",
                 116,
                 
                 P
                 , 
                 
                 35520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011011; B = 8'b11111100; // Expected: {'P': 55188}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011011; B = 8'b11111100; | Outputs: P=%b | Expected: P=%d",
                 117,
                 
                 P
                 , 
                 
                 55188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010111; B = 8'b10100011; // Expected: {'P': 14181}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010111; B = 8'b10100011; | Outputs: P=%b | Expected: P=%d",
                 118,
                 
                 P
                 , 
                 
                 14181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100010; B = 8'b10011101; // Expected: {'P': 5338}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100010; B = 8'b10011101; | Outputs: P=%b | Expected: P=%d",
                 119,
                 
                 P
                 , 
                 
                 5338
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111110; B = 8'b11111101; // Expected: {'P': 15686}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111110; B = 8'b11111101; | Outputs: P=%b | Expected: P=%d",
                 120,
                 
                 P
                 , 
                 
                 15686
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100000; B = 8'b11010011; // Expected: {'P': 33760}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100000; B = 8'b11010011; | Outputs: P=%b | Expected: P=%d",
                 121,
                 
                 P
                 , 
                 
                 33760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000000; B = 8'b00111111; // Expected: {'P': 8064}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000000; B = 8'b00111111; | Outputs: P=%b | Expected: P=%d",
                 122,
                 
                 P
                 , 
                 
                 8064
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100101; B = 8'b11111100; // Expected: {'P': 41580}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100101; B = 8'b11111100; | Outputs: P=%b | Expected: P=%d",
                 123,
                 
                 P
                 , 
                 
                 41580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000000; B = 8'b00111101; // Expected: {'P': 11712}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000000; B = 8'b00111101; | Outputs: P=%b | Expected: P=%d",
                 124,
                 
                 P
                 , 
                 
                 11712
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001011; B = 8'b00110111; // Expected: {'P': 605}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001011; B = 8'b00110111; | Outputs: P=%b | Expected: P=%d",
                 125,
                 
                 P
                 , 
                 
                 605
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110101; B = 8'b10101011; // Expected: {'P': 41895}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110101; B = 8'b10101011; | Outputs: P=%b | Expected: P=%d",
                 126,
                 
                 P
                 , 
                 
                 41895
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011010; B = 8'b10101101; // Expected: {'P': 26642}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011010; B = 8'b10101101; | Outputs: P=%b | Expected: P=%d",
                 127,
                 
                 P
                 , 
                 
                 26642
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101011; B = 8'b10010110; // Expected: {'P': 25650}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101011; B = 8'b10010110; | Outputs: P=%b | Expected: P=%d",
                 128,
                 
                 P
                 , 
                 
                 25650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100011; B = 8'b10111110; // Expected: {'P': 6650}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100011; B = 8'b10111110; | Outputs: P=%b | Expected: P=%d",
                 129,
                 
                 P
                 , 
                 
                 6650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000110; B = 8'b00010110; // Expected: {'P': 2948}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000110; B = 8'b00010110; | Outputs: P=%b | Expected: P=%d",
                 130,
                 
                 P
                 , 
                 
                 2948
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110000; B = 8'b10101010; // Expected: {'P': 29920}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110000; B = 8'b10101010; | Outputs: P=%b | Expected: P=%d",
                 131,
                 
                 P
                 , 
                 
                 29920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110001; B = 8'b01010010; // Expected: {'P': 4018}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110001; B = 8'b01010010; | Outputs: P=%b | Expected: P=%d",
                 132,
                 
                 P
                 , 
                 
                 4018
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010001; B = 8'b00011000; // Expected: {'P': 408}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010001; B = 8'b00011000; | Outputs: P=%b | Expected: P=%d",
                 133,
                 
                 P
                 , 
                 
                 408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101100; B = 8'b10101001; // Expected: {'P': 7436}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101100; B = 8'b10101001; | Outputs: P=%b | Expected: P=%d",
                 134,
                 
                 P
                 , 
                 
                 7436
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000001; B = 8'b10111011; // Expected: {'P': 36091}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000001; B = 8'b10111011; | Outputs: P=%b | Expected: P=%d",
                 135,
                 
                 P
                 , 
                 
                 36091
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101011; B = 8'b11010010; // Expected: {'P': 49350}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101011; B = 8'b11010010; | Outputs: P=%b | Expected: P=%d",
                 136,
                 
                 P
                 , 
                 
                 49350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011011; B = 8'b11110010; // Expected: {'P': 6534}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011011; B = 8'b11110010; | Outputs: P=%b | Expected: P=%d",
                 137,
                 
                 P
                 , 
                 
                 6534
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101110; B = 8'b11000101; // Expected: {'P': 21670}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101110; B = 8'b11000101; | Outputs: P=%b | Expected: P=%d",
                 138,
                 
                 P
                 , 
                 
                 21670
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001101; B = 8'b10010000; // Expected: {'P': 1872}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001101; B = 8'b10010000; | Outputs: P=%b | Expected: P=%d",
                 139,
                 
                 P
                 , 
                 
                 1872
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101111; B = 8'b11110001; // Expected: {'P': 57599}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101111; B = 8'b11110001; | Outputs: P=%b | Expected: P=%d",
                 140,
                 
                 P
                 , 
                 
                 57599
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010100; B = 8'b01010101; // Expected: {'P': 1700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010100; B = 8'b01010101; | Outputs: P=%b | Expected: P=%d",
                 141,
                 
                 P
                 , 
                 
                 1700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101111; B = 8'b10010100; // Expected: {'P': 16428}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101111; B = 8'b10010100; | Outputs: P=%b | Expected: P=%d",
                 142,
                 
                 P
                 , 
                 
                 16428
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110001; B = 8'b11111011; // Expected: {'P': 60491}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110001; B = 8'b11111011; | Outputs: P=%b | Expected: P=%d",
                 143,
                 
                 P
                 , 
                 
                 60491
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111100; B = 8'b10111101; // Expected: {'P': 47628}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111100; B = 8'b10111101; | Outputs: P=%b | Expected: P=%d",
                 144,
                 
                 P
                 , 
                 
                 47628
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000110; B = 8'b10010111; // Expected: {'P': 10570}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000110; B = 8'b10010111; | Outputs: P=%b | Expected: P=%d",
                 145,
                 
                 P
                 , 
                 
                 10570
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010101; B = 8'b00101011; // Expected: {'P': 9159}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010101; B = 8'b00101011; | Outputs: P=%b | Expected: P=%d",
                 146,
                 
                 P
                 , 
                 
                 9159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011101; B = 8'b11110000; // Expected: {'P': 37680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011101; B = 8'b11110000; | Outputs: P=%b | Expected: P=%d",
                 147,
                 
                 P
                 , 
                 
                 37680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111111; B = 8'b01010101; // Expected: {'P': 21675}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111111; B = 8'b01010101; | Outputs: P=%b | Expected: P=%d",
                 148,
                 
                 P
                 , 
                 
                 21675
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111010; B = 8'b11110010; // Expected: {'P': 60500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111010; B = 8'b11110010; | Outputs: P=%b | Expected: P=%d",
                 149,
                 
                 P
                 , 
                 
                 60500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010001; B = 8'b11100010; // Expected: {'P': 47234}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010001; B = 8'b11100010; | Outputs: P=%b | Expected: P=%d",
                 150,
                 
                 P
                 , 
                 
                 47234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111100; B = 8'b01101010; // Expected: {'P': 6360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111100; B = 8'b01101010; | Outputs: P=%b | Expected: P=%d",
                 151,
                 
                 P
                 , 
                 
                 6360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111101; B = 8'b11100110; // Expected: {'P': 28750}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111101; B = 8'b11100110; | Outputs: P=%b | Expected: P=%d",
                 152,
                 
                 P
                 , 
                 
                 28750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011111; B = 8'b11011101; // Expected: {'P': 49283}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011111; B = 8'b11011101; | Outputs: P=%b | Expected: P=%d",
                 153,
                 
                 P
                 , 
                 
                 49283
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100110; B = 8'b01101000; // Expected: {'P': 17264}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100110; B = 8'b01101000; | Outputs: P=%b | Expected: P=%d",
                 154,
                 
                 P
                 , 
                 
                 17264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110010; B = 8'b11000100; // Expected: {'P': 34888}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110010; B = 8'b11000100; | Outputs: P=%b | Expected: P=%d",
                 155,
                 
                 P
                 , 
                 
                 34888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011111; B = 8'b01001011; // Expected: {'P': 11925}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011111; B = 8'b01001011; | Outputs: P=%b | Expected: P=%d",
                 156,
                 
                 P
                 , 
                 
                 11925
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011001; B = 8'b10010100; // Expected: {'P': 32116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011001; B = 8'b10010100; | Outputs: P=%b | Expected: P=%d",
                 157,
                 
                 P
                 , 
                 
                 32116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111010; B = 8'b10000001; // Expected: {'P': 23994}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111010; B = 8'b10000001; | Outputs: P=%b | Expected: P=%d",
                 158,
                 
                 P
                 , 
                 
                 23994
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111011; B = 8'b11011011; // Expected: {'P': 26937}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111011; B = 8'b11011011; | Outputs: P=%b | Expected: P=%d",
                 159,
                 
                 P
                 , 
                 
                 26937
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000001; B = 8'b00011110; // Expected: {'P': 1950}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000001; B = 8'b00011110; | Outputs: P=%b | Expected: P=%d",
                 160,
                 
                 P
                 , 
                 
                 1950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101101; B = 8'b10010011; // Expected: {'P': 6615}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101101; B = 8'b10010011; | Outputs: P=%b | Expected: P=%d",
                 161,
                 
                 P
                 , 
                 
                 6615
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111000; B = 8'b11010100; // Expected: {'P': 52576}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111000; B = 8'b11010100; | Outputs: P=%b | Expected: P=%d",
                 162,
                 
                 P
                 , 
                 
                 52576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101100; B = 8'b01011010; // Expected: {'P': 3960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101100; B = 8'b01011010; | Outputs: P=%b | Expected: P=%d",
                 163,
                 
                 P
                 , 
                 
                 3960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010100; B = 8'b10010011; // Expected: {'P': 21756}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010100; B = 8'b10010011; | Outputs: P=%b | Expected: P=%d",
                 164,
                 
                 P
                 , 
                 
                 21756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100100; B = 8'b10010010; // Expected: {'P': 14600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100100; B = 8'b10010010; | Outputs: P=%b | Expected: P=%d",
                 165,
                 
                 P
                 , 
                 
                 14600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000011; B = 8'b11110111; // Expected: {'P': 32357}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000011; B = 8'b11110111; | Outputs: P=%b | Expected: P=%d",
                 166,
                 
                 P
                 , 
                 
                 32357
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010111; B = 8'b10011000; // Expected: {'P': 13224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010111; B = 8'b10011000; | Outputs: P=%b | Expected: P=%d",
                 167,
                 
                 P
                 , 
                 
                 13224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111111; B = 8'b01100010; // Expected: {'P': 18718}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111111; B = 8'b01100010; | Outputs: P=%b | Expected: P=%d",
                 168,
                 
                 P
                 , 
                 
                 18718
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100000; B = 8'b00101110; // Expected: {'P': 4416}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100000; B = 8'b00101110; | Outputs: P=%b | Expected: P=%d",
                 169,
                 
                 P
                 , 
                 
                 4416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000001; B = 8'b11001000; // Expected: {'P': 38600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000001; B = 8'b11001000; | Outputs: P=%b | Expected: P=%d",
                 170,
                 
                 P
                 , 
                 
                 38600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000001; B = 8'b11011011; // Expected: {'P': 219}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000001; B = 8'b11011011; | Outputs: P=%b | Expected: P=%d",
                 171,
                 
                 P
                 , 
                 
                 219
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100001; B = 8'b10011001; // Expected: {'P': 5049}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100001; B = 8'b10011001; | Outputs: P=%b | Expected: P=%d",
                 172,
                 
                 P
                 , 
                 
                 5049
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000010; B = 8'b10000011; // Expected: {'P': 262}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000010; B = 8'b10000011; | Outputs: P=%b | Expected: P=%d",
                 173,
                 
                 P
                 , 
                 
                 262
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010011; B = 8'b10111000; // Expected: {'P': 15272}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010011; B = 8'b10111000; | Outputs: P=%b | Expected: P=%d",
                 174,
                 
                 P
                 , 
                 
                 15272
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100011; B = 8'b00000101; // Expected: {'P': 175}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100011; B = 8'b00000101; | Outputs: P=%b | Expected: P=%d",
                 175,
                 
                 P
                 , 
                 
                 175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100111; B = 8'b10011110; // Expected: {'P': 26386}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100111; B = 8'b10011110; | Outputs: P=%b | Expected: P=%d",
                 176,
                 
                 P
                 , 
                 
                 26386
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111100; B = 8'b11100010; // Expected: {'P': 42488}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111100; B = 8'b11100010; | Outputs: P=%b | Expected: P=%d",
                 177,
                 
                 P
                 , 
                 
                 42488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001111; B = 8'b11101111; // Expected: {'P': 3585}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001111; B = 8'b11101111; | Outputs: P=%b | Expected: P=%d",
                 178,
                 
                 P
                 , 
                 
                 3585
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110010; B = 8'b00110001; // Expected: {'P': 8722}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110010; B = 8'b00110001; | Outputs: P=%b | Expected: P=%d",
                 179,
                 
                 P
                 , 
                 
                 8722
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011010; B = 8'b00000101; // Expected: {'P': 450}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011010; B = 8'b00000101; | Outputs: P=%b | Expected: P=%d",
                 180,
                 
                 P
                 , 
                 
                 450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010111; B = 8'b01000100; // Expected: {'P': 5916}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010111; B = 8'b01000100; | Outputs: P=%b | Expected: P=%d",
                 181,
                 
                 P
                 , 
                 
                 5916
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100001; B = 8'b11010010; // Expected: {'P': 47250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100001; B = 8'b11010010; | Outputs: P=%b | Expected: P=%d",
                 182,
                 
                 P
                 , 
                 
                 47250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001101; B = 8'b11010110; // Expected: {'P': 30174}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001101; B = 8'b11010110; | Outputs: P=%b | Expected: P=%d",
                 183,
                 
                 P
                 , 
                 
                 30174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001010; B = 8'b11111000; // Expected: {'P': 34224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001010; B = 8'b11111000; | Outputs: P=%b | Expected: P=%d",
                 184,
                 
                 P
                 , 
                 
                 34224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100001; B = 8'b11011100; // Expected: {'P': 35420}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100001; B = 8'b11011100; | Outputs: P=%b | Expected: P=%d",
                 185,
                 
                 P
                 , 
                 
                 35420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110010; B = 8'b10101101; // Expected: {'P': 30794}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110010; B = 8'b10101101; | Outputs: P=%b | Expected: P=%d",
                 186,
                 
                 P
                 , 
                 
                 30794
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001010; B = 8'b10111110; // Expected: {'P': 26220}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001010; B = 8'b10111110; | Outputs: P=%b | Expected: P=%d",
                 187,
                 
                 P
                 , 
                 
                 26220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010111; B = 8'b01101110; // Expected: {'P': 16610}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010111; B = 8'b01101110; | Outputs: P=%b | Expected: P=%d",
                 188,
                 
                 P
                 , 
                 
                 16610
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010101; B = 8'b11101110; // Expected: {'P': 50694}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010101; B = 8'b11101110; | Outputs: P=%b | Expected: P=%d",
                 189,
                 
                 P
                 , 
                 
                 50694
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111111; B = 8'b00000001; // Expected: {'P': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111111; B = 8'b00000001; | Outputs: P=%b | Expected: P=%d",
                 190,
                 
                 P
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110111; B = 8'b11101000; // Expected: {'P': 12760}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110111; B = 8'b11101000; | Outputs: P=%b | Expected: P=%d",
                 191,
                 
                 P
                 , 
                 
                 12760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010000; B = 8'b10101100; // Expected: {'P': 13760}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010000; B = 8'b10101100; | Outputs: P=%b | Expected: P=%d",
                 192,
                 
                 P
                 , 
                 
                 13760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011110; B = 8'b10111111; // Expected: {'P': 17954}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011110; B = 8'b10111111; | Outputs: P=%b | Expected: P=%d",
                 193,
                 
                 P
                 , 
                 
                 17954
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000101; B = 8'b10110010; // Expected: {'P': 12282}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000101; B = 8'b10110010; | Outputs: P=%b | Expected: P=%d",
                 194,
                 
                 P
                 , 
                 
                 12282
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001100; B = 8'b11010111; // Expected: {'P': 2580}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001100; B = 8'b11010111; | Outputs: P=%b | Expected: P=%d",
                 195,
                 
                 P
                 , 
                 
                 2580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001111; B = 8'b01101000; // Expected: {'P': 14872}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001111; B = 8'b01101000; | Outputs: P=%b | Expected: P=%d",
                 196,
                 
                 P
                 , 
                 
                 14872
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010101; B = 8'b01000101; // Expected: {'P': 5865}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010101; B = 8'b01000101; | Outputs: P=%b | Expected: P=%d",
                 197,
                 
                 P
                 , 
                 
                 5865
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101101; B = 8'b00001110; // Expected: {'P': 3318}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101101; B = 8'b00001110; | Outputs: P=%b | Expected: P=%d",
                 198,
                 
                 P
                 , 
                 
                 3318
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101111; B = 8'b00011101; // Expected: {'P': 1363}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101111; B = 8'b00011101; | Outputs: P=%b | Expected: P=%d",
                 199,
                 
                 P
                 , 
                 
                 1363
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101101; B = 8'b01011100; // Expected: {'P': 4140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101101; B = 8'b01011100; | Outputs: P=%b | Expected: P=%d",
                 200,
                 
                 P
                 , 
                 
                 4140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100010; B = 8'b10111000; // Expected: {'P': 41584}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100010; B = 8'b10111000; | Outputs: P=%b | Expected: P=%d",
                 201,
                 
                 P
                 , 
                 
                 41584
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111011; B = 8'b11010111; // Expected: {'P': 26445}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111011; B = 8'b11010111; | Outputs: P=%b | Expected: P=%d",
                 202,
                 
                 P
                 , 
                 
                 26445
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000111; B = 8'b01101011; // Expected: {'P': 749}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000111; B = 8'b01101011; | Outputs: P=%b | Expected: P=%d",
                 203,
                 
                 P
                 , 
                 
                 749
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101000; B = 8'b10001110; // Expected: {'P': 5680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101000; B = 8'b10001110; | Outputs: P=%b | Expected: P=%d",
                 204,
                 
                 P
                 , 
                 
                 5680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001010; B = 8'b00000100; // Expected: {'P': 808}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001010; B = 8'b00000100; | Outputs: P=%b | Expected: P=%d",
                 205,
                 
                 P
                 , 
                 
                 808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101010; B = 8'b00010101; // Expected: {'P': 4914}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101010; B = 8'b00010101; | Outputs: P=%b | Expected: P=%d",
                 206,
                 
                 P
                 , 
                 
                 4914
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101001; B = 8'b01111000; // Expected: {'P': 12600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101001; B = 8'b01111000; | Outputs: P=%b | Expected: P=%d",
                 207,
                 
                 P
                 , 
                 
                 12600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010001; B = 8'b10010011; // Expected: {'P': 30723}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010001; B = 8'b10010011; | Outputs: P=%b | Expected: P=%d",
                 208,
                 
                 P
                 , 
                 
                 30723
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001000; B = 8'b01001111; // Expected: {'P': 15800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001000; B = 8'b01001111; | Outputs: P=%b | Expected: P=%d",
                 209,
                 
                 P
                 , 
                 
                 15800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000101; B = 8'b00100011; // Expected: {'P': 4655}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000101; B = 8'b00100011; | Outputs: P=%b | Expected: P=%d",
                 210,
                 
                 P
                 , 
                 
                 4655
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000100; B = 8'b01010001; // Expected: {'P': 15876}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000100; B = 8'b01010001; | Outputs: P=%b | Expected: P=%d",
                 211,
                 
                 P
                 , 
                 
                 15876
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011111; B = 8'b01000001; // Expected: {'P': 14495}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011111; B = 8'b01000001; | Outputs: P=%b | Expected: P=%d",
                 212,
                 
                 P
                 , 
                 
                 14495
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111111; B = 8'b10000101; // Expected: {'P': 8379}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111111; B = 8'b10000101; | Outputs: P=%b | Expected: P=%d",
                 213,
                 
                 P
                 , 
                 
                 8379
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101011; B = 8'b01000000; // Expected: {'P': 6848}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101011; B = 8'b01000000; | Outputs: P=%b | Expected: P=%d",
                 214,
                 
                 P
                 , 
                 
                 6848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101100; B = 8'b10001101; // Expected: {'P': 6204}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101100; B = 8'b10001101; | Outputs: P=%b | Expected: P=%d",
                 215,
                 
                 P
                 , 
                 
                 6204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110011; B = 8'b00100010; // Expected: {'P': 8262}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110011; B = 8'b00100010; | Outputs: P=%b | Expected: P=%d",
                 216,
                 
                 P
                 , 
                 
                 8262
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000001; B = 8'b00101111; // Expected: {'P': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000001; B = 8'b00101111; | Outputs: P=%b | Expected: P=%d",
                 217,
                 
                 P
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110001; B = 8'b01001111; // Expected: {'P': 19039}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110001; B = 8'b01001111; | Outputs: P=%b | Expected: P=%d",
                 218,
                 
                 P
                 , 
                 
                 19039
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001001; B = 8'b11101010; // Expected: {'P': 47034}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001001; B = 8'b11101010; | Outputs: P=%b | Expected: P=%d",
                 219,
                 
                 P
                 , 
                 
                 47034
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101111; B = 8'b00010010; // Expected: {'P': 4302}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101111; B = 8'b00010010; | Outputs: P=%b | Expected: P=%d",
                 220,
                 
                 P
                 , 
                 
                 4302
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010001; B = 8'b11000001; // Expected: {'P': 15633}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010001; B = 8'b11000001; | Outputs: P=%b | Expected: P=%d",
                 221,
                 
                 P
                 , 
                 
                 15633
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001100; B = 8'b11010111; // Expected: {'P': 43860}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001100; B = 8'b11010111; | Outputs: P=%b | Expected: P=%d",
                 222,
                 
                 P
                 , 
                 
                 43860
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110011; B = 8'b01011111; // Expected: {'P': 10925}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110011; B = 8'b01011111; | Outputs: P=%b | Expected: P=%d",
                 223,
                 
                 P
                 , 
                 
                 10925
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000011; B = 8'b11001001; // Expected: {'P': 26331}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000011; B = 8'b11001001; | Outputs: P=%b | Expected: P=%d",
                 224,
                 
                 P
                 , 
                 
                 26331
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100110; B = 8'b01010111; // Expected: {'P': 3306}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100110; B = 8'b01010111; | Outputs: P=%b | Expected: P=%d",
                 225,
                 
                 P
                 , 
                 
                 3306
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011010; B = 8'b00101010; // Expected: {'P': 6468}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011010; B = 8'b00101010; | Outputs: P=%b | Expected: P=%d",
                 226,
                 
                 P
                 , 
                 
                 6468
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000110; B = 8'b11100001; // Expected: {'P': 30150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000110; B = 8'b11100001; | Outputs: P=%b | Expected: P=%d",
                 227,
                 
                 P
                 , 
                 
                 30150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010100; B = 8'b01000011; // Expected: {'P': 14204}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010100; B = 8'b01000011; | Outputs: P=%b | Expected: P=%d",
                 228,
                 
                 P
                 , 
                 
                 14204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100000; B = 8'b01010010; // Expected: {'P': 13120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100000; B = 8'b01010010; | Outputs: P=%b | Expected: P=%d",
                 229,
                 
                 P
                 , 
                 
                 13120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010100; B = 8'b10001110; // Expected: {'P': 2840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010100; B = 8'b10001110; | Outputs: P=%b | Expected: P=%d",
                 230,
                 
                 P
                 , 
                 
                 2840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000111; B = 8'b10100101; // Expected: {'P': 32835}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000111; B = 8'b10100101; | Outputs: P=%b | Expected: P=%d",
                 231,
                 
                 P
                 , 
                 
                 32835
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100001; B = 8'b11110000; // Expected: {'P': 7920}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100001; B = 8'b11110000; | Outputs: P=%b | Expected: P=%d",
                 232,
                 
                 P
                 , 
                 
                 7920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111011; B = 8'b10001011; // Expected: {'P': 34889}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111011; B = 8'b10001011; | Outputs: P=%b | Expected: P=%d",
                 233,
                 
                 P
                 , 
                 
                 34889
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100011; B = 8'b01100111; // Expected: {'P': 10197}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100011; B = 8'b01100111; | Outputs: P=%b | Expected: P=%d",
                 234,
                 
                 P
                 , 
                 
                 10197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011011; B = 8'b01111000; // Expected: {'P': 18600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011011; B = 8'b01111000; | Outputs: P=%b | Expected: P=%d",
                 235,
                 
                 P
                 , 
                 
                 18600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111010; B = 8'b00110000; // Expected: {'P': 2784}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111010; B = 8'b00110000; | Outputs: P=%b | Expected: P=%d",
                 236,
                 
                 P
                 , 
                 
                 2784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100011; B = 8'b00010011; // Expected: {'P': 665}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100011; B = 8'b00010011; | Outputs: P=%b | Expected: P=%d",
                 237,
                 
                 P
                 , 
                 
                 665
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100010; B = 8'b10000010; // Expected: {'P': 4420}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100010; B = 8'b10000010; | Outputs: P=%b | Expected: P=%d",
                 238,
                 
                 P
                 , 
                 
                 4420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111111; B = 8'b11000111; // Expected: {'P': 50745}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111111; B = 8'b11000111; | Outputs: P=%b | Expected: P=%d",
                 239,
                 
                 P
                 , 
                 
                 50745
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110101; B = 8'b11001011; // Expected: {'P': 23751}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110101; B = 8'b11001011; | Outputs: P=%b | Expected: P=%d",
                 240,
                 
                 P
                 , 
                 
                 23751
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000101; B = 8'b01001100; // Expected: {'P': 5244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000101; B = 8'b01001100; | Outputs: P=%b | Expected: P=%d",
                 241,
                 
                 P
                 , 
                 
                 5244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011010; B = 8'b11000011; // Expected: {'P': 5070}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011010; B = 8'b11000011; | Outputs: P=%b | Expected: P=%d",
                 242,
                 
                 P
                 , 
                 
                 5070
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011010; B = 8'b11111010; // Expected: {'P': 22500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011010; B = 8'b11111010; | Outputs: P=%b | Expected: P=%d",
                 243,
                 
                 P
                 , 
                 
                 22500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000011; B = 8'b00010100; // Expected: {'P': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000011; B = 8'b00010100; | Outputs: P=%b | Expected: P=%d",
                 244,
                 
                 P
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100000; B = 8'b10001101; // Expected: {'P': 22560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100000; B = 8'b10001101; | Outputs: P=%b | Expected: P=%d",
                 245,
                 
                 P
                 , 
                 
                 22560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111101; B = 8'b01000111; // Expected: {'P': 4331}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111101; B = 8'b01000111; | Outputs: P=%b | Expected: P=%d",
                 246,
                 
                 P
                 , 
                 
                 4331
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100001; B = 8'b10010100; // Expected: {'P': 14356}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100001; B = 8'b10010100; | Outputs: P=%b | Expected: P=%d",
                 247,
                 
                 P
                 , 
                 
                 14356
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111101; B = 8'b01001111; // Expected: {'P': 4819}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111101; B = 8'b01001111; | Outputs: P=%b | Expected: P=%d",
                 248,
                 
                 P
                 , 
                 
                 4819
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011111; B = 8'b01111001; // Expected: {'P': 26983}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011111; B = 8'b01111001; | Outputs: P=%b | Expected: P=%d",
                 249,
                 
                 P
                 , 
                 
                 26983
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001110; B = 8'b00011111; // Expected: {'P': 4402}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001110; B = 8'b00011111; | Outputs: P=%b | Expected: P=%d",
                 250,
                 
                 P
                 , 
                 
                 4402
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101101; B = 8'b00111100; // Expected: {'P': 14220}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101101; B = 8'b00111100; | Outputs: P=%b | Expected: P=%d",
                 251,
                 
                 P
                 , 
                 
                 14220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101100; B = 8'b11010001; // Expected: {'P': 49324}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101100; B = 8'b11010001; | Outputs: P=%b | Expected: P=%d",
                 252,
                 
                 P
                 , 
                 
                 49324
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011000; B = 8'b11010100; // Expected: {'P': 32224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011000; B = 8'b11010100; | Outputs: P=%b | Expected: P=%d",
                 253,
                 
                 P
                 , 
                 
                 32224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100000; B = 8'b01101110; // Expected: {'P': 24640}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100000; B = 8'b01101110; | Outputs: P=%b | Expected: P=%d",
                 254,
                 
                 P
                 , 
                 
                 24640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110110; B = 8'b00110010; // Expected: {'P': 9100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110110; B = 8'b00110010; | Outputs: P=%b | Expected: P=%d",
                 255,
                 
                 P
                 , 
                 
                 9100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100001; B = 8'b01000101; // Expected: {'P': 2277}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100001; B = 8'b01000101; | Outputs: P=%b | Expected: P=%d",
                 256,
                 
                 P
                 , 
                 
                 2277
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110100; B = 8'b11101010; // Expected: {'P': 12168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110100; B = 8'b11101010; | Outputs: P=%b | Expected: P=%d",
                 257,
                 
                 P
                 , 
                 
                 12168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011001; B = 8'b01011110; // Expected: {'P': 14382}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011001; B = 8'b01011110; | Outputs: P=%b | Expected: P=%d",
                 258,
                 
                 P
                 , 
                 
                 14382
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001001; B = 8'b00000111; // Expected: {'P': 959}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001001; B = 8'b00000111; | Outputs: P=%b | Expected: P=%d",
                 259,
                 
                 P
                 , 
                 
                 959
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000101; B = 8'b11000001; // Expected: {'P': 965}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000101; B = 8'b11000001; | Outputs: P=%b | Expected: P=%d",
                 260,
                 
                 P
                 , 
                 
                 965
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010111; B = 8'b01110010; // Expected: {'P': 24510}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010111; B = 8'b01110010; | Outputs: P=%b | Expected: P=%d",
                 261,
                 
                 P
                 , 
                 
                 24510
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001111; B = 8'b11011100; // Expected: {'P': 45540}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001111; B = 8'b11011100; | Outputs: P=%b | Expected: P=%d",
                 262,
                 
                 P
                 , 
                 
                 45540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111010; B = 8'b11011001; // Expected: {'P': 40362}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111010; B = 8'b11011001; | Outputs: P=%b | Expected: P=%d",
                 263,
                 
                 P
                 , 
                 
                 40362
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111000; B = 8'b11010101; // Expected: {'P': 39192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111000; B = 8'b11010101; | Outputs: P=%b | Expected: P=%d",
                 264,
                 
                 P
                 , 
                 
                 39192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001100; B = 8'b11111011; // Expected: {'P': 35140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001100; B = 8'b11111011; | Outputs: P=%b | Expected: P=%d",
                 265,
                 
                 P
                 , 
                 
                 35140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100000; B = 8'b00011011; // Expected: {'P': 2592}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100000; B = 8'b00011011; | Outputs: P=%b | Expected: P=%d",
                 266,
                 
                 P
                 , 
                 
                 2592
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010000; B = 8'b11110100; // Expected: {'P': 19520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010000; B = 8'b11110100; | Outputs: P=%b | Expected: P=%d",
                 267,
                 
                 P
                 , 
                 
                 19520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110111; B = 8'b01011000; // Expected: {'P': 10472}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110111; B = 8'b01011000; | Outputs: P=%b | Expected: P=%d",
                 268,
                 
                 P
                 , 
                 
                 10472
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111111; B = 8'b11000010; // Expected: {'P': 49470}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111111; B = 8'b11000010; | Outputs: P=%b | Expected: P=%d",
                 269,
                 
                 P
                 , 
                 
                 49470
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011100; B = 8'b00110110; // Expected: {'P': 1512}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011100; B = 8'b00110110; | Outputs: P=%b | Expected: P=%d",
                 270,
                 
                 P
                 , 
                 
                 1512
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111001; B = 8'b00010011; // Expected: {'P': 3515}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111001; B = 8'b00010011; | Outputs: P=%b | Expected: P=%d",
                 271,
                 
                 P
                 , 
                 
                 3515
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101000; B = 8'b00000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101000; B = 8'b00000000; | Outputs: P=%b | Expected: P=%d",
                 272,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110100; B = 8'b01100100; // Expected: {'P': 11600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110100; B = 8'b01100100; | Outputs: P=%b | Expected: P=%d",
                 273,
                 
                 P
                 , 
                 
                 11600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100010; B = 8'b01100001; // Expected: {'P': 9506}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100010; B = 8'b01100001; | Outputs: P=%b | Expected: P=%d",
                 274,
                 
                 P
                 , 
                 
                 9506
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111110; B = 8'b10110100; // Expected: {'P': 45720}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111110; B = 8'b10110100; | Outputs: P=%b | Expected: P=%d",
                 275,
                 
                 P
                 , 
                 
                 45720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101101; B = 8'b11001011; // Expected: {'P': 22127}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101101; B = 8'b11001011; | Outputs: P=%b | Expected: P=%d",
                 276,
                 
                 P
                 , 
                 
                 22127
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101101; B = 8'b01011011; // Expected: {'P': 15743}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101101; B = 8'b01011011; | Outputs: P=%b | Expected: P=%d",
                 277,
                 
                 P
                 , 
                 
                 15743
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110010; B = 8'b11110001; // Expected: {'P': 58322}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110010; B = 8'b11110001; | Outputs: P=%b | Expected: P=%d",
                 278,
                 
                 P
                 , 
                 
                 58322
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100010; B = 8'b11011011; // Expected: {'P': 35478}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100010; B = 8'b11011011; | Outputs: P=%b | Expected: P=%d",
                 279,
                 
                 P
                 , 
                 
                 35478
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111000; B = 8'b01110110; // Expected: {'P': 21712}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111000; B = 8'b01110110; | Outputs: P=%b | Expected: P=%d",
                 280,
                 
                 P
                 , 
                 
                 21712
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111101; B = 8'b01110111; // Expected: {'P': 22491}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111101; B = 8'b01110111; | Outputs: P=%b | Expected: P=%d",
                 281,
                 
                 P
                 , 
                 
                 22491
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011111; B = 8'b11111010; // Expected: {'P': 7750}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011111; B = 8'b11111010; | Outputs: P=%b | Expected: P=%d",
                 282,
                 
                 P
                 , 
                 
                 7750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100111; B = 8'b01011011; // Expected: {'P': 3549}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100111; B = 8'b01011011; | Outputs: P=%b | Expected: P=%d",
                 283,
                 
                 P
                 , 
                 
                 3549
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000110; B = 8'b11000001; // Expected: {'P': 38214}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000110; B = 8'b11000001; | Outputs: P=%b | Expected: P=%d",
                 284,
                 
                 P
                 , 
                 
                 38214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110111; B = 8'b01011110; // Expected: {'P': 17202}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110111; B = 8'b01011110; | Outputs: P=%b | Expected: P=%d",
                 285,
                 
                 P
                 , 
                 
                 17202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111001; B = 8'b11001010; // Expected: {'P': 24442}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111001; B = 8'b11001010; | Outputs: P=%b | Expected: P=%d",
                 286,
                 
                 P
                 , 
                 
                 24442
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010011; B = 8'b01101000; // Expected: {'P': 8632}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010011; B = 8'b01101000; | Outputs: P=%b | Expected: P=%d",
                 287,
                 
                 P
                 , 
                 
                 8632
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011011; B = 8'b10010000; // Expected: {'P': 3888}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011011; B = 8'b10010000; | Outputs: P=%b | Expected: P=%d",
                 288,
                 
                 P
                 , 
                 
                 3888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101110; B = 8'b11001010; // Expected: {'P': 48076}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101110; B = 8'b11001010; | Outputs: P=%b | Expected: P=%d",
                 289,
                 
                 P
                 , 
                 
                 48076
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100011; B = 8'b01011001; // Expected: {'P': 8811}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100011; B = 8'b01011001; | Outputs: P=%b | Expected: P=%d",
                 290,
                 
                 P
                 , 
                 
                 8811
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011001; B = 8'b11100011; // Expected: {'P': 49259}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011001; B = 8'b11100011; | Outputs: P=%b | Expected: P=%d",
                 291,
                 
                 P
                 , 
                 
                 49259
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011010; B = 8'b00000010; // Expected: {'P': 308}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011010; B = 8'b00000010; | Outputs: P=%b | Expected: P=%d",
                 292,
                 
                 P
                 , 
                 
                 308
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011001; B = 8'b11000011; // Expected: {'P': 42315}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011001; B = 8'b11000011; | Outputs: P=%b | Expected: P=%d",
                 293,
                 
                 P
                 , 
                 
                 42315
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001110; B = 8'b11011000; // Expected: {'P': 16848}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001110; B = 8'b11011000; | Outputs: P=%b | Expected: P=%d",
                 294,
                 
                 P
                 , 
                 
                 16848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100010; B = 8'b00011100; // Expected: {'P': 6328}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100010; B = 8'b00011100; | Outputs: P=%b | Expected: P=%d",
                 295,
                 
                 P
                 , 
                 
                 6328
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001100; B = 8'b00011111; // Expected: {'P': 372}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001100; B = 8'b00011111; | Outputs: P=%b | Expected: P=%d",
                 296,
                 
                 P
                 , 
                 
                 372
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100001; B = 8'b00100010; // Expected: {'P': 1122}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100001; B = 8'b00100010; | Outputs: P=%b | Expected: P=%d",
                 297,
                 
                 P
                 , 
                 
                 1122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110100; B = 8'b11011011; // Expected: {'P': 39420}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110100; B = 8'b11011011; | Outputs: P=%b | Expected: P=%d",
                 298,
                 
                 P
                 , 
                 
                 39420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101011; B = 8'b11100000; // Expected: {'P': 23968}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101011; B = 8'b11100000; | Outputs: P=%b | Expected: P=%d",
                 299,
                 
                 P
                 , 
                 
                 23968
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000011; B = 8'b11011110; // Expected: {'P': 666}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000011; B = 8'b11011110; | Outputs: P=%b | Expected: P=%d",
                 300,
                 
                 P
                 , 
                 
                 666
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000101; B = 8'b10100000; // Expected: {'P': 800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000101; B = 8'b10100000; | Outputs: P=%b | Expected: P=%d",
                 301,
                 
                 P
                 , 
                 
                 800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101000; B = 8'b01101000; // Expected: {'P': 10816}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101000; B = 8'b01101000; | Outputs: P=%b | Expected: P=%d",
                 302,
                 
                 P
                 , 
                 
                 10816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001000; B = 8'b10001000; // Expected: {'P': 27200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001000; B = 8'b10001000; | Outputs: P=%b | Expected: P=%d",
                 303,
                 
                 P
                 , 
                 
                 27200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101111; B = 8'b01111101; // Expected: {'P': 29875}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101111; B = 8'b01111101; | Outputs: P=%b | Expected: P=%d",
                 304,
                 
                 P
                 , 
                 
                 29875
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010010; B = 8'b01111111; // Expected: {'P': 2286}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010010; B = 8'b01111111; | Outputs: P=%b | Expected: P=%d",
                 305,
                 
                 P
                 , 
                 
                 2286
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010100; B = 8'b10100101; // Expected: {'P': 13860}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010100; B = 8'b10100101; | Outputs: P=%b | Expected: P=%d",
                 306,
                 
                 P
                 , 
                 
                 13860
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011000; B = 8'b00110110; // Expected: {'P': 11664}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011000; B = 8'b00110110; | Outputs: P=%b | Expected: P=%d",
                 307,
                 
                 P
                 , 
                 
                 11664
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101011; B = 8'b10010100; // Expected: {'P': 6364}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101011; B = 8'b10010100; | Outputs: P=%b | Expected: P=%d",
                 308,
                 
                 P
                 , 
                 
                 6364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001110; B = 8'b00100110; // Expected: {'P': 7828}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001110; B = 8'b00100110; | Outputs: P=%b | Expected: P=%d",
                 309,
                 
                 P
                 , 
                 
                 7828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010100; B = 8'b00111010; // Expected: {'P': 12296}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010100; B = 8'b00111010; | Outputs: P=%b | Expected: P=%d",
                 310,
                 
                 P
                 , 
                 
                 12296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010001; B = 8'b11011001; // Expected: {'P': 45353}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010001; B = 8'b11011001; | Outputs: P=%b | Expected: P=%d",
                 311,
                 
                 P
                 , 
                 
                 45353
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110101; B = 8'b00100111; // Expected: {'P': 4563}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110101; B = 8'b00100111; | Outputs: P=%b | Expected: P=%d",
                 312,
                 
                 P
                 , 
                 
                 4563
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101000; B = 8'b11010101; // Expected: {'P': 35784}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101000; B = 8'b11010101; | Outputs: P=%b | Expected: P=%d",
                 313,
                 
                 P
                 , 
                 
                 35784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011010; B = 8'b10110010; // Expected: {'P': 27412}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011010; B = 8'b10110010; | Outputs: P=%b | Expected: P=%d",
                 314,
                 
                 P
                 , 
                 
                 27412
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001001; B = 8'b11100111; // Expected: {'P': 16863}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001001; B = 8'b11100111; | Outputs: P=%b | Expected: P=%d",
                 315,
                 
                 P
                 , 
                 
                 16863
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101101; B = 8'b10011000; // Expected: {'P': 16568}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101101; B = 8'b10011000; | Outputs: P=%b | Expected: P=%d",
                 316,
                 
                 P
                 , 
                 
                 16568
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110110; B = 8'b01111010; // Expected: {'P': 14396}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110110; B = 8'b01111010; | Outputs: P=%b | Expected: P=%d",
                 317,
                 
                 P
                 , 
                 
                 14396
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010100; B = 8'b10101111; // Expected: {'P': 37100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010100; B = 8'b10101111; | Outputs: P=%b | Expected: P=%d",
                 318,
                 
                 P
                 , 
                 
                 37100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101110; B = 8'b01100001; // Expected: {'P': 10670}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101110; B = 8'b01100001; | Outputs: P=%b | Expected: P=%d",
                 319,
                 
                 P
                 , 
                 
                 10670
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001001; B = 8'b01100110; // Expected: {'P': 918}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001001; B = 8'b01100110; | Outputs: P=%b | Expected: P=%d",
                 320,
                 
                 P
                 , 
                 
                 918
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110001; B = 8'b11000110; // Expected: {'P': 47718}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110001; B = 8'b11000110; | Outputs: P=%b | Expected: P=%d",
                 321,
                 
                 P
                 , 
                 
                 47718
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101111; B = 8'b01000101; // Expected: {'P': 3243}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101111; B = 8'b01000101; | Outputs: P=%b | Expected: P=%d",
                 322,
                 
                 P
                 , 
                 
                 3243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000001; B = 8'b01100111; // Expected: {'P': 103}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000001; B = 8'b01100111; | Outputs: P=%b | Expected: P=%d",
                 323,
                 
                 P
                 , 
                 
                 103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001100; B = 8'b00101010; // Expected: {'P': 8568}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001100; B = 8'b00101010; | Outputs: P=%b | Expected: P=%d",
                 324,
                 
                 P
                 , 
                 
                 8568
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111011; B = 8'b00011110; // Expected: {'P': 5610}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111011; B = 8'b00011110; | Outputs: P=%b | Expected: P=%d",
                 325,
                 
                 P
                 , 
                 
                 5610
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110101; B = 8'b00101001; // Expected: {'P': 10045}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110101; B = 8'b00101001; | Outputs: P=%b | Expected: P=%d",
                 326,
                 
                 P
                 , 
                 
                 10045
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111010; B = 8'b11100111; // Expected: {'P': 57750}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111010; B = 8'b11100111; | Outputs: P=%b | Expected: P=%d",
                 327,
                 
                 P
                 , 
                 
                 57750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111001; B = 8'b10010110; // Expected: {'P': 37350}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111001; B = 8'b10010110; | Outputs: P=%b | Expected: P=%d",
                 328,
                 
                 P
                 , 
                 
                 37350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111010; B = 8'b01010011; // Expected: {'P': 4814}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111010; B = 8'b01010011; | Outputs: P=%b | Expected: P=%d",
                 329,
                 
                 P
                 , 
                 
                 4814
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001111; B = 8'b00011111; // Expected: {'P': 465}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001111; B = 8'b00011111; | Outputs: P=%b | Expected: P=%d",
                 330,
                 
                 P
                 , 
                 
                 465
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010010; B = 8'b01100110; // Expected: {'P': 1836}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010010; B = 8'b01100110; | Outputs: P=%b | Expected: P=%d",
                 331,
                 
                 P
                 , 
                 
                 1836
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010000; B = 8'b00000011; // Expected: {'P': 432}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010000; B = 8'b00000011; | Outputs: P=%b | Expected: P=%d",
                 332,
                 
                 P
                 , 
                 
                 432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111010; B = 8'b01111100; // Expected: {'P': 7192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111010; B = 8'b01111100; | Outputs: P=%b | Expected: P=%d",
                 333,
                 
                 P
                 , 
                 
                 7192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010111; B = 8'b00000110; // Expected: {'P': 906}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010111; B = 8'b00000110; | Outputs: P=%b | Expected: P=%d",
                 334,
                 
                 P
                 , 
                 
                 906
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101111; B = 8'b11111100; // Expected: {'P': 44100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101111; B = 8'b11111100; | Outputs: P=%b | Expected: P=%d",
                 335,
                 
                 P
                 , 
                 
                 44100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011010; B = 8'b01010100; // Expected: {'P': 7560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011010; B = 8'b01010100; | Outputs: P=%b | Expected: P=%d",
                 336,
                 
                 P
                 , 
                 
                 7560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000000; B = 8'b10100100; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000000; B = 8'b10100100; | Outputs: P=%b | Expected: P=%d",
                 337,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010010; B = 8'b10110000; // Expected: {'P': 36960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010010; B = 8'b10110000; | Outputs: P=%b | Expected: P=%d",
                 338,
                 
                 P
                 , 
                 
                 36960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011111; B = 8'b11011000; // Expected: {'P': 34344}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011111; B = 8'b11011000; | Outputs: P=%b | Expected: P=%d",
                 339,
                 
                 P
                 , 
                 
                 34344
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010000; B = 8'b00100111; // Expected: {'P': 8112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010000; B = 8'b00100111; | Outputs: P=%b | Expected: P=%d",
                 340,
                 
                 P
                 , 
                 
                 8112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011010; B = 8'b11001100; // Expected: {'P': 31416}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011010; B = 8'b11001100; | Outputs: P=%b | Expected: P=%d",
                 341,
                 
                 P
                 , 
                 
                 31416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110110; B = 8'b00110001; // Expected: {'P': 12054}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110110; B = 8'b00110001; | Outputs: P=%b | Expected: P=%d",
                 342,
                 
                 P
                 , 
                 
                 12054
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110001; B = 8'b11110010; // Expected: {'P': 11858}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110001; B = 8'b11110010; | Outputs: P=%b | Expected: P=%d",
                 343,
                 
                 P
                 , 
                 
                 11858
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011010; B = 8'b01000010; // Expected: {'P': 5940}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011010; B = 8'b01000010; | Outputs: P=%b | Expected: P=%d",
                 344,
                 
                 P
                 , 
                 
                 5940
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101000; B = 8'b10111000; // Expected: {'P': 7360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101000; B = 8'b10111000; | Outputs: P=%b | Expected: P=%d",
                 345,
                 
                 P
                 , 
                 
                 7360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001011; B = 8'b11101010; // Expected: {'P': 47502}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001011; B = 8'b11101010; | Outputs: P=%b | Expected: P=%d",
                 346,
                 
                 P
                 , 
                 
                 47502
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000001; B = 8'b01001101; // Expected: {'P': 14861}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000001; B = 8'b01001101; | Outputs: P=%b | Expected: P=%d",
                 347,
                 
                 P
                 , 
                 
                 14861
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111000; B = 8'b10101001; // Expected: {'P': 9464}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111000; B = 8'b10101001; | Outputs: P=%b | Expected: P=%d",
                 348,
                 
                 P
                 , 
                 
                 9464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000011; B = 8'b01010110; // Expected: {'P': 16770}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000011; B = 8'b01010110; | Outputs: P=%b | Expected: P=%d",
                 349,
                 
                 P
                 , 
                 
                 16770
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001000; B = 8'b01100000; // Expected: {'P': 6912}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001000; B = 8'b01100000; | Outputs: P=%b | Expected: P=%d",
                 350,
                 
                 P
                 , 
                 
                 6912
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110101; B = 8'b10110010; // Expected: {'P': 20826}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110101; B = 8'b10110010; | Outputs: P=%b | Expected: P=%d",
                 351,
                 
                 P
                 , 
                 
                 20826
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100100; B = 8'b00110110; // Expected: {'P': 12312}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100100; B = 8'b00110110; | Outputs: P=%b | Expected: P=%d",
                 352,
                 
                 P
                 , 
                 
                 12312
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011100; B = 8'b10001010; // Expected: {'P': 12696}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011100; B = 8'b10001010; | Outputs: P=%b | Expected: P=%d",
                 353,
                 
                 P
                 , 
                 
                 12696
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111101; B = 8'b01100000; // Expected: {'P': 24288}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111101; B = 8'b01100000; | Outputs: P=%b | Expected: P=%d",
                 354,
                 
                 P
                 , 
                 
                 24288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011100; B = 8'b10000110; // Expected: {'P': 3752}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011100; B = 8'b10000110; | Outputs: P=%b | Expected: P=%d",
                 355,
                 
                 P
                 , 
                 
                 3752
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010110; B = 8'b10010110; // Expected: {'P': 32100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010110; B = 8'b10010110; | Outputs: P=%b | Expected: P=%d",
                 356,
                 
                 P
                 , 
                 
                 32100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111000; B = 8'b00010000; // Expected: {'P': 896}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111000; B = 8'b00010000; | Outputs: P=%b | Expected: P=%d",
                 357,
                 
                 P
                 , 
                 
                 896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000101; B = 8'b10100001; // Expected: {'P': 11109}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000101; B = 8'b10100001; | Outputs: P=%b | Expected: P=%d",
                 358,
                 
                 P
                 , 
                 
                 11109
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010110; B = 8'b00111010; // Expected: {'P': 4988}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010110; B = 8'b00111010; | Outputs: P=%b | Expected: P=%d",
                 359,
                 
                 P
                 , 
                 
                 4988
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110101; B = 8'b10010101; // Expected: {'P': 26969}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110101; B = 8'b10010101; | Outputs: P=%b | Expected: P=%d",
                 360,
                 
                 P
                 , 
                 
                 26969
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000010; B = 8'b01100100; // Expected: {'P': 19400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000010; B = 8'b01100100; | Outputs: P=%b | Expected: P=%d",
                 361,
                 
                 P
                 , 
                 
                 19400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111100; B = 8'b00000011; // Expected: {'P': 564}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111100; B = 8'b00000011; | Outputs: P=%b | Expected: P=%d",
                 362,
                 
                 P
                 , 
                 
                 564
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001110; B = 8'b00010001; // Expected: {'P': 238}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001110; B = 8'b00010001; | Outputs: P=%b | Expected: P=%d",
                 363,
                 
                 P
                 , 
                 
                 238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011110; B = 8'b10000011; // Expected: {'P': 12314}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011110; B = 8'b10000011; | Outputs: P=%b | Expected: P=%d",
                 364,
                 
                 P
                 , 
                 
                 12314
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100111; B = 8'b00001110; // Expected: {'P': 1442}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100111; B = 8'b00001110; | Outputs: P=%b | Expected: P=%d",
                 365,
                 
                 P
                 , 
                 
                 1442
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110101; B = 8'b00011001; // Expected: {'P': 6125}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110101; B = 8'b00011001; | Outputs: P=%b | Expected: P=%d",
                 366,
                 
                 P
                 , 
                 
                 6125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111110; B = 8'b11110011; // Expected: {'P': 15066}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111110; B = 8'b11110011; | Outputs: P=%b | Expected: P=%d",
                 367,
                 
                 P
                 , 
                 
                 15066
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100100; B = 8'b01110001; // Expected: {'P': 18532}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100100; B = 8'b01110001; | Outputs: P=%b | Expected: P=%d",
                 368,
                 
                 P
                 , 
                 
                 18532
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100011; B = 8'b11100100; // Expected: {'P': 7980}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100011; B = 8'b11100100; | Outputs: P=%b | Expected: P=%d",
                 369,
                 
                 P
                 , 
                 
                 7980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000100; B = 8'b01010100; // Expected: {'P': 16464}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000100; B = 8'b01010100; | Outputs: P=%b | Expected: P=%d",
                 370,
                 
                 P
                 , 
                 
                 16464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110110; B = 8'b10110101; // Expected: {'P': 32942}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110110; B = 8'b10110101; | Outputs: P=%b | Expected: P=%d",
                 371,
                 
                 P
                 , 
                 
                 32942
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000010; B = 8'b00001110; // Expected: {'P': 2716}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000010; B = 8'b00001110; | Outputs: P=%b | Expected: P=%d",
                 372,
                 
                 P
                 , 
                 
                 2716
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011001; B = 8'b01010000; // Expected: {'P': 7120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011001; B = 8'b01010000; | Outputs: P=%b | Expected: P=%d",
                 373,
                 
                 P
                 , 
                 
                 7120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001000; B = 8'b11001110; // Expected: {'P': 28016}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001000; B = 8'b11001110; | Outputs: P=%b | Expected: P=%d",
                 374,
                 
                 P
                 , 
                 
                 28016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011000; B = 8'b00001011; // Expected: {'P': 968}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011000; B = 8'b00001011; | Outputs: P=%b | Expected: P=%d",
                 375,
                 
                 P
                 , 
                 
                 968
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110011; B = 8'b10000110; // Expected: {'P': 15410}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110011; B = 8'b10000110; | Outputs: P=%b | Expected: P=%d",
                 376,
                 
                 P
                 , 
                 
                 15410
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001000; B = 8'b11000111; // Expected: {'P': 1592}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001000; B = 8'b11000111; | Outputs: P=%b | Expected: P=%d",
                 377,
                 
                 P
                 , 
                 
                 1592
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110110; B = 8'b00101001; // Expected: {'P': 2214}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110110; B = 8'b00101001; | Outputs: P=%b | Expected: P=%d",
                 378,
                 
                 P
                 , 
                 
                 2214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111011; B = 8'b11101101; // Expected: {'P': 13983}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111011; B = 8'b11101101; | Outputs: P=%b | Expected: P=%d",
                 379,
                 
                 P
                 , 
                 
                 13983
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111001; B = 8'b11000011; // Expected: {'P': 23595}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111001; B = 8'b11000011; | Outputs: P=%b | Expected: P=%d",
                 380,
                 
                 P
                 , 
                 
                 23595
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001001; B = 8'b10011111; // Expected: {'P': 1431}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001001; B = 8'b10011111; | Outputs: P=%b | Expected: P=%d",
                 381,
                 
                 P
                 , 
                 
                 1431
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100110; B = 8'b00110111; // Expected: {'P': 12650}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100110; B = 8'b00110111; | Outputs: P=%b | Expected: P=%d",
                 382,
                 
                 P
                 , 
                 
                 12650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011001; B = 8'b01101010; // Expected: {'P': 16218}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011001; B = 8'b01101010; | Outputs: P=%b | Expected: P=%d",
                 383,
                 
                 P
                 , 
                 
                 16218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100110; B = 8'b01110110; // Expected: {'P': 4484}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100110; B = 8'b01110110; | Outputs: P=%b | Expected: P=%d",
                 384,
                 
                 P
                 , 
                 
                 4484
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001100; B = 8'b01100110; // Expected: {'P': 7752}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001100; B = 8'b01100110; | Outputs: P=%b | Expected: P=%d",
                 385,
                 
                 P
                 , 
                 
                 7752
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100100; B = 8'b01001010; // Expected: {'P': 7400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100100; B = 8'b01001010; | Outputs: P=%b | Expected: P=%d",
                 386,
                 
                 P
                 , 
                 
                 7400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001101; B = 8'b00100110; // Expected: {'P': 5358}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001101; B = 8'b00100110; | Outputs: P=%b | Expected: P=%d",
                 387,
                 
                 P
                 , 
                 
                 5358
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000110; B = 8'b01110110; // Expected: {'P': 23364}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000110; B = 8'b01110110; | Outputs: P=%b | Expected: P=%d",
                 388,
                 
                 P
                 , 
                 
                 23364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110100; B = 8'b00101111; // Expected: {'P': 11468}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110100; B = 8'b00101111; | Outputs: P=%b | Expected: P=%d",
                 389,
                 
                 P
                 , 
                 
                 11468
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110010; B = 8'b01001001; // Expected: {'P': 8322}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110010; B = 8'b01001001; | Outputs: P=%b | Expected: P=%d",
                 390,
                 
                 P
                 , 
                 
                 8322
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000001; B = 8'b00011110; // Expected: {'P': 5790}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000001; B = 8'b00011110; | Outputs: P=%b | Expected: P=%d",
                 391,
                 
                 P
                 , 
                 
                 5790
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001000; B = 8'b10000000; // Expected: {'P': 17408}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001000; B = 8'b10000000; | Outputs: P=%b | Expected: P=%d",
                 392,
                 
                 P
                 , 
                 
                 17408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001110; B = 8'b00111001; // Expected: {'P': 798}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001110; B = 8'b00111001; | Outputs: P=%b | Expected: P=%d",
                 393,
                 
                 P
                 , 
                 
                 798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010100; B = 8'b11101000; // Expected: {'P': 4640}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010100; B = 8'b11101000; | Outputs: P=%b | Expected: P=%d",
                 394,
                 
                 P
                 , 
                 
                 4640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011100; B = 8'b00110001; // Expected: {'P': 7644}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011100; B = 8'b00110001; | Outputs: P=%b | Expected: P=%d",
                 395,
                 
                 P
                 , 
                 
                 7644
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011100; B = 8'b11110011; // Expected: {'P': 6804}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011100; B = 8'b11110011; | Outputs: P=%b | Expected: P=%d",
                 396,
                 
                 P
                 , 
                 
                 6804
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010110; B = 8'b00001101; // Expected: {'P': 1950}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010110; B = 8'b00001101; | Outputs: P=%b | Expected: P=%d",
                 397,
                 
                 P
                 , 
                 
                 1950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100110; B = 8'b01101001; // Expected: {'P': 17430}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100110; B = 8'b01101001; | Outputs: P=%b | Expected: P=%d",
                 398,
                 
                 P
                 , 
                 
                 17430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100111; B = 8'b10011111; // Expected: {'P': 16377}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100111; B = 8'b10011111; | Outputs: P=%b | Expected: P=%d",
                 399,
                 
                 P
                 , 
                 
                 16377
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100100; B = 8'b11011110; // Expected: {'P': 7992}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100100; B = 8'b11011110; | Outputs: P=%b | Expected: P=%d",
                 400,
                 
                 P
                 , 
                 
                 7992
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011010; B = 8'b01100010; // Expected: {'P': 15092}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011010; B = 8'b01100010; | Outputs: P=%b | Expected: P=%d",
                 401,
                 
                 P
                 , 
                 
                 15092
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110011; B = 8'b01011101; // Expected: {'P': 16647}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110011; B = 8'b01011101; | Outputs: P=%b | Expected: P=%d",
                 402,
                 
                 P
                 , 
                 
                 16647
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111000; B = 8'b01100111; // Expected: {'P': 5768}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111000; B = 8'b01100111; | Outputs: P=%b | Expected: P=%d",
                 403,
                 
                 P
                 , 
                 
                 5768
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000101; B = 8'b00100000; // Expected: {'P': 4256}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000101; B = 8'b00100000; | Outputs: P=%b | Expected: P=%d",
                 404,
                 
                 P
                 , 
                 
                 4256
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000110; B = 8'b11100000; // Expected: {'P': 30016}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000110; B = 8'b11100000; | Outputs: P=%b | Expected: P=%d",
                 405,
                 
                 P
                 , 
                 
                 30016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001100; B = 8'b11101010; // Expected: {'P': 32760}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001100; B = 8'b11101010; | Outputs: P=%b | Expected: P=%d",
                 406,
                 
                 P
                 , 
                 
                 32760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010010; B = 8'b11110011; // Expected: {'P': 35478}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010010; B = 8'b11110011; | Outputs: P=%b | Expected: P=%d",
                 407,
                 
                 P
                 , 
                 
                 35478
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000111; B = 8'b11111001; // Expected: {'P': 17679}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000111; B = 8'b11111001; | Outputs: P=%b | Expected: P=%d",
                 408,
                 
                 P
                 , 
                 
                 17679
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010111; B = 8'b01010011; // Expected: {'P': 7221}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010111; B = 8'b01010011; | Outputs: P=%b | Expected: P=%d",
                 409,
                 
                 P
                 , 
                 
                 7221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101011; B = 8'b00101000; // Expected: {'P': 1720}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101011; B = 8'b00101000; | Outputs: P=%b | Expected: P=%d",
                 410,
                 
                 P
                 , 
                 
                 1720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110010; B = 8'b11011011; // Expected: {'P': 10950}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110010; B = 8'b11011011; | Outputs: P=%b | Expected: P=%d",
                 411,
                 
                 P
                 , 
                 
                 10950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101100; B = 8'b10100100; // Expected: {'P': 17712}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101100; B = 8'b10100100; | Outputs: P=%b | Expected: P=%d",
                 412,
                 
                 P
                 , 
                 
                 17712
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000011; B = 8'b10111010; // Expected: {'P': 24366}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000011; B = 8'b10111010; | Outputs: P=%b | Expected: P=%d",
                 413,
                 
                 P
                 , 
                 
                 24366
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000111; B = 8'b01010010; // Expected: {'P': 5822}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000111; B = 8'b01010010; | Outputs: P=%b | Expected: P=%d",
                 414,
                 
                 P
                 , 
                 
                 5822
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101110; B = 8'b01100010; // Expected: {'P': 10780}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101110; B = 8'b01100010; | Outputs: P=%b | Expected: P=%d",
                 415,
                 
                 P
                 , 
                 
                 10780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111010; B = 8'b01110011; // Expected: {'P': 6670}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111010; B = 8'b01110011; | Outputs: P=%b | Expected: P=%d",
                 416,
                 
                 P
                 , 
                 
                 6670
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110111; B = 8'b00110111; // Expected: {'P': 10065}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110111; B = 8'b00110111; | Outputs: P=%b | Expected: P=%d",
                 417,
                 
                 P
                 , 
                 
                 10065
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111001; B = 8'b01000010; // Expected: {'P': 16434}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111001; B = 8'b01000010; | Outputs: P=%b | Expected: P=%d",
                 418,
                 
                 P
                 , 
                 
                 16434
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110010; B = 8'b10111010; // Expected: {'P': 45012}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110010; B = 8'b10111010; | Outputs: P=%b | Expected: P=%d",
                 419,
                 
                 P
                 , 
                 
                 45012
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110010; B = 8'b01000000; // Expected: {'P': 11392}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110010; B = 8'b01000000; | Outputs: P=%b | Expected: P=%d",
                 420,
                 
                 P
                 , 
                 
                 11392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000010; B = 8'b00011100; // Expected: {'P': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000010; B = 8'b00011100; | Outputs: P=%b | Expected: P=%d",
                 421,
                 
                 P
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110100; B = 8'b11000110; // Expected: {'P': 22968}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110100; B = 8'b11000110; | Outputs: P=%b | Expected: P=%d",
                 422,
                 
                 P
                 , 
                 
                 22968
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110000; B = 8'b01110110; // Expected: {'P': 13216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110000; B = 8'b01110110; | Outputs: P=%b | Expected: P=%d",
                 423,
                 
                 P
                 , 
                 
                 13216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101111; B = 8'b01000000; // Expected: {'P': 15296}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101111; B = 8'b01000000; | Outputs: P=%b | Expected: P=%d",
                 424,
                 
                 P
                 , 
                 
                 15296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110111; B = 8'b10011011; // Expected: {'P': 8525}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110111; B = 8'b10011011; | Outputs: P=%b | Expected: P=%d",
                 425,
                 
                 P
                 , 
                 
                 8525
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111100; B = 8'b10110010; // Expected: {'P': 33464}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111100; B = 8'b10110010; | Outputs: P=%b | Expected: P=%d",
                 426,
                 
                 P
                 , 
                 
                 33464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101000; B = 8'b00001000; // Expected: {'P': 1856}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101000; B = 8'b00001000; | Outputs: P=%b | Expected: P=%d",
                 427,
                 
                 P
                 , 
                 
                 1856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011111; B = 8'b11010001; // Expected: {'P': 33231}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011111; B = 8'b11010001; | Outputs: P=%b | Expected: P=%d",
                 428,
                 
                 P
                 , 
                 
                 33231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100100; B = 8'b11010100; // Expected: {'P': 48336}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100100; B = 8'b11010100; | Outputs: P=%b | Expected: P=%d",
                 429,
                 
                 P
                 , 
                 
                 48336
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100010; B = 8'b10110100; // Expected: {'P': 40680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100010; B = 8'b10110100; | Outputs: P=%b | Expected: P=%d",
                 430,
                 
                 P
                 , 
                 
                 40680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011100; B = 8'b11010110; // Expected: {'P': 5992}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011100; B = 8'b11010110; | Outputs: P=%b | Expected: P=%d",
                 431,
                 
                 P
                 , 
                 
                 5992
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110101; B = 8'b11101011; // Expected: {'P': 27495}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110101; B = 8'b11101011; | Outputs: P=%b | Expected: P=%d",
                 432,
                 
                 P
                 , 
                 
                 27495
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100011; B = 8'b01000101; // Expected: {'P': 2415}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100011; B = 8'b01000101; | Outputs: P=%b | Expected: P=%d",
                 433,
                 
                 P
                 , 
                 
                 2415
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100000; B = 8'b01011001; // Expected: {'P': 2848}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100000; B = 8'b01011001; | Outputs: P=%b | Expected: P=%d",
                 434,
                 
                 P
                 , 
                 
                 2848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101010; B = 8'b00111110; // Expected: {'P': 2604}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101010; B = 8'b00111110; | Outputs: P=%b | Expected: P=%d",
                 435,
                 
                 P
                 , 
                 
                 2604
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000000; B = 8'b01001100; // Expected: {'P': 9728}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000000; B = 8'b01001100; | Outputs: P=%b | Expected: P=%d",
                 436,
                 
                 P
                 , 
                 
                 9728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101001; B = 8'b01010100; // Expected: {'P': 3444}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101001; B = 8'b01010100; | Outputs: P=%b | Expected: P=%d",
                 437,
                 
                 P
                 , 
                 
                 3444
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100100; B = 8'b10101000; // Expected: {'P': 6048}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100100; B = 8'b10101000; | Outputs: P=%b | Expected: P=%d",
                 438,
                 
                 P
                 , 
                 
                 6048
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011110; B = 8'b00100101; // Expected: {'P': 5846}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011110; B = 8'b00100101; | Outputs: P=%b | Expected: P=%d",
                 439,
                 
                 P
                 , 
                 
                 5846
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111111; B = 8'b00110010; // Expected: {'P': 3150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111111; B = 8'b00110010; | Outputs: P=%b | Expected: P=%d",
                 440,
                 
                 P
                 , 
                 
                 3150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100111; B = 8'b11000111; // Expected: {'P': 33233}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100111; B = 8'b11000111; | Outputs: P=%b | Expected: P=%d",
                 441,
                 
                 P
                 , 
                 
                 33233
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001010; B = 8'b01011010; // Expected: {'P': 900}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001010; B = 8'b01011010; | Outputs: P=%b | Expected: P=%d",
                 442,
                 
                 P
                 , 
                 
                 900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101100; B = 8'b10001100; // Expected: {'P': 24080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101100; B = 8'b10001100; | Outputs: P=%b | Expected: P=%d",
                 443,
                 
                 P
                 , 
                 
                 24080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101111; B = 8'b11110000; // Expected: {'P': 42000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101111; B = 8'b11110000; | Outputs: P=%b | Expected: P=%d",
                 444,
                 
                 P
                 , 
                 
                 42000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100010; B = 8'b00000100; // Expected: {'P': 648}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100010; B = 8'b00000100; | Outputs: P=%b | Expected: P=%d",
                 445,
                 
                 P
                 , 
                 
                 648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011110; B = 8'b11000010; // Expected: {'P': 30652}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011110; B = 8'b11000010; | Outputs: P=%b | Expected: P=%d",
                 446,
                 
                 P
                 , 
                 
                 30652
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100100; B = 8'b10010000; // Expected: {'P': 23616}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100100; B = 8'b10010000; | Outputs: P=%b | Expected: P=%d",
                 447,
                 
                 P
                 , 
                 
                 23616
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000101; B = 8'b01011111; // Expected: {'P': 6555}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000101; B = 8'b01011111; | Outputs: P=%b | Expected: P=%d",
                 448,
                 
                 P
                 , 
                 
                 6555
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101010; B = 8'b10101111; // Expected: {'P': 18550}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101010; B = 8'b10101111; | Outputs: P=%b | Expected: P=%d",
                 449,
                 
                 P
                 , 
                 
                 18550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000101; B = 8'b01101101; // Expected: {'P': 14497}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000101; B = 8'b01101101; | Outputs: P=%b | Expected: P=%d",
                 450,
                 
                 P
                 , 
                 
                 14497
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000111; B = 8'b10111100; // Expected: {'P': 25380}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000111; B = 8'b10111100; | Outputs: P=%b | Expected: P=%d",
                 451,
                 
                 P
                 , 
                 
                 25380
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010101; B = 8'b00010110; // Expected: {'P': 4686}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010101; B = 8'b00010110; | Outputs: P=%b | Expected: P=%d",
                 452,
                 
                 P
                 , 
                 
                 4686
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001010; B = 8'b00010100; // Expected: {'P': 1480}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001010; B = 8'b00010100; | Outputs: P=%b | Expected: P=%d",
                 453,
                 
                 P
                 , 
                 
                 1480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010001; B = 8'b11001101; // Expected: {'P': 42845}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010001; B = 8'b11001101; | Outputs: P=%b | Expected: P=%d",
                 454,
                 
                 P
                 , 
                 
                 42845
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011011; B = 8'b10000101; // Expected: {'P': 3591}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011011; B = 8'b10000101; | Outputs: P=%b | Expected: P=%d",
                 455,
                 
                 P
                 , 
                 
                 3591
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110010; B = 8'b00001101; // Expected: {'P': 2314}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110010; B = 8'b00001101; | Outputs: P=%b | Expected: P=%d",
                 456,
                 
                 P
                 , 
                 
                 2314
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100000; B = 8'b10110011; // Expected: {'P': 5728}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100000; B = 8'b10110011; | Outputs: P=%b | Expected: P=%d",
                 457,
                 
                 P
                 , 
                 
                 5728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110111; B = 8'b11101110; // Expected: {'P': 58786}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110111; B = 8'b11101110; | Outputs: P=%b | Expected: P=%d",
                 458,
                 
                 P
                 , 
                 
                 58786
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101001; B = 8'b01011111; // Expected: {'P': 3895}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101001; B = 8'b01011111; | Outputs: P=%b | Expected: P=%d",
                 459,
                 
                 P
                 , 
                 
                 3895
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000001; B = 8'b01100110; // Expected: {'P': 19686}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000001; B = 8'b01100110; | Outputs: P=%b | Expected: P=%d",
                 460,
                 
                 P
                 , 
                 
                 19686
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011111; B = 8'b11110010; // Expected: {'P': 7502}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011111; B = 8'b11110010; | Outputs: P=%b | Expected: P=%d",
                 461,
                 
                 P
                 , 
                 
                 7502
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011111; B = 8'b00100000; // Expected: {'P': 3040}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011111; B = 8'b00100000; | Outputs: P=%b | Expected: P=%d",
                 462,
                 
                 P
                 , 
                 
                 3040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110000; B = 8'b01111010; // Expected: {'P': 5856}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110000; B = 8'b01111010; | Outputs: P=%b | Expected: P=%d",
                 463,
                 
                 P
                 , 
                 
                 5856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011111; B = 8'b10101001; // Expected: {'P': 16055}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011111; B = 8'b10101001; | Outputs: P=%b | Expected: P=%d",
                 464,
                 
                 P
                 , 
                 
                 16055
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001001; B = 8'b01110010; // Expected: {'P': 22914}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001001; B = 8'b01110010; | Outputs: P=%b | Expected: P=%d",
                 465,
                 
                 P
                 , 
                 
                 22914
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110001; B = 8'b01101111; // Expected: {'P': 12543}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110001; B = 8'b01101111; | Outputs: P=%b | Expected: P=%d",
                 466,
                 
                 P
                 , 
                 
                 12543
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001000; B = 8'b10010000; // Expected: {'P': 28800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001000; B = 8'b10010000; | Outputs: P=%b | Expected: P=%d",
                 467,
                 
                 P
                 , 
                 
                 28800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111111; B = 8'b10100011; // Expected: {'P': 31133}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111111; B = 8'b10100011; | Outputs: P=%b | Expected: P=%d",
                 468,
                 
                 P
                 , 
                 
                 31133
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111101; B = 8'b00101100; // Expected: {'P': 8316}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111101; B = 8'b00101100; | Outputs: P=%b | Expected: P=%d",
                 469,
                 
                 P
                 , 
                 
                 8316
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110101; B = 8'b00011000; // Expected: {'P': 1272}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110101; B = 8'b00011000; | Outputs: P=%b | Expected: P=%d",
                 470,
                 
                 P
                 , 
                 
                 1272
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001000; B = 8'b10011011; // Expected: {'P': 11160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001000; B = 8'b10011011; | Outputs: P=%b | Expected: P=%d",
                 471,
                 
                 P
                 , 
                 
                 11160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111010; B = 8'b10001000; // Expected: {'P': 7888}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111010; B = 8'b10001000; | Outputs: P=%b | Expected: P=%d",
                 472,
                 
                 P
                 , 
                 
                 7888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001101; B = 8'b11001001; // Expected: {'P': 28341}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001101; B = 8'b11001001; | Outputs: P=%b | Expected: P=%d",
                 473,
                 
                 P
                 , 
                 
                 28341
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010011; B = 8'b01100101; // Expected: {'P': 1919}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010011; B = 8'b01100101; | Outputs: P=%b | Expected: P=%d",
                 474,
                 
                 P
                 , 
                 
                 1919
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010100; B = 8'b11001101; // Expected: {'P': 30340}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010100; B = 8'b11001101; | Outputs: P=%b | Expected: P=%d",
                 475,
                 
                 P
                 , 
                 
                 30340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101101; B = 8'b11011111; // Expected: {'P': 24307}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101101; B = 8'b11011111; | Outputs: P=%b | Expected: P=%d",
                 476,
                 
                 P
                 , 
                 
                 24307
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011110; B = 8'b10100101; // Expected: {'P': 26070}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011110; B = 8'b10100101; | Outputs: P=%b | Expected: P=%d",
                 477,
                 
                 P
                 , 
                 
                 26070
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101000; B = 8'b00001010; // Expected: {'P': 1680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101000; B = 8'b00001010; | Outputs: P=%b | Expected: P=%d",
                 478,
                 
                 P
                 , 
                 
                 1680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100001; B = 8'b01011001; // Expected: {'P': 20025}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100001; B = 8'b01011001; | Outputs: P=%b | Expected: P=%d",
                 479,
                 
                 P
                 , 
                 
                 20025
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100110; B = 8'b10110111; // Expected: {'P': 30378}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100110; B = 8'b10110111; | Outputs: P=%b | Expected: P=%d",
                 480,
                 
                 P
                 , 
                 
                 30378
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100011; B = 8'b00111111; // Expected: {'P': 10269}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100011; B = 8'b00111111; | Outputs: P=%b | Expected: P=%d",
                 481,
                 
                 P
                 , 
                 
                 10269
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100001; B = 8'b00111110; // Expected: {'P': 9982}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100001; B = 8'b00111110; | Outputs: P=%b | Expected: P=%d",
                 482,
                 
                 P
                 , 
                 
                 9982
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000011; B = 8'b01000010; // Expected: {'P': 12870}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000011; B = 8'b01000010; | Outputs: P=%b | Expected: P=%d",
                 483,
                 
                 P
                 , 
                 
                 12870
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100111; B = 8'b10100000; // Expected: {'P': 6240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100111; B = 8'b10100000; | Outputs: P=%b | Expected: P=%d",
                 484,
                 
                 P
                 , 
                 
                 6240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111100; B = 8'b10010011; // Expected: {'P': 37044}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111100; B = 8'b10010011; | Outputs: P=%b | Expected: P=%d",
                 485,
                 
                 P
                 , 
                 
                 37044
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101100; B = 8'b10101011; // Expected: {'P': 18468}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101100; B = 8'b10101011; | Outputs: P=%b | Expected: P=%d",
                 486,
                 
                 P
                 , 
                 
                 18468
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100000; B = 8'b01000100; // Expected: {'P': 15232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100000; B = 8'b01000100; | Outputs: P=%b | Expected: P=%d",
                 487,
                 
                 P
                 , 
                 
                 15232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010010; B = 8'b10010101; // Expected: {'P': 21754}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010010; B = 8'b10010101; | Outputs: P=%b | Expected: P=%d",
                 488,
                 
                 P
                 , 
                 
                 21754
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011010; B = 8'b01101000; // Expected: {'P': 16016}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011010; B = 8'b01101000; | Outputs: P=%b | Expected: P=%d",
                 489,
                 
                 P
                 , 
                 
                 16016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011111; B = 8'b01111010; // Expected: {'P': 3782}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011111; B = 8'b01111010; | Outputs: P=%b | Expected: P=%d",
                 490,
                 
                 P
                 , 
                 
                 3782
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110101; B = 8'b00111100; // Expected: {'P': 10860}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110101; B = 8'b00111100; | Outputs: P=%b | Expected: P=%d",
                 491,
                 
                 P
                 , 
                 
                 10860
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011101; B = 8'b00100001; // Expected: {'P': 5181}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011101; B = 8'b00100001; | Outputs: P=%b | Expected: P=%d",
                 492,
                 
                 P
                 , 
                 
                 5181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011001; B = 8'b11111000; // Expected: {'P': 37944}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011001; B = 8'b11111000; | Outputs: P=%b | Expected: P=%d",
                 493,
                 
                 P
                 , 
                 
                 37944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100011; B = 8'b00100100; // Expected: {'P': 8172}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100011; B = 8'b00100100; | Outputs: P=%b | Expected: P=%d",
                 494,
                 
                 P
                 , 
                 
                 8172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101100; B = 8'b01011110; // Expected: {'P': 10152}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101100; B = 8'b01011110; | Outputs: P=%b | Expected: P=%d",
                 495,
                 
                 P
                 , 
                 
                 10152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010111; B = 8'b00001101; // Expected: {'P': 2795}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010111; B = 8'b00001101; | Outputs: P=%b | Expected: P=%d",
                 496,
                 
                 P
                 , 
                 
                 2795
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000101; B = 8'b01110110; // Expected: {'P': 23246}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000101; B = 8'b01110110; | Outputs: P=%b | Expected: P=%d",
                 497,
                 
                 P
                 , 
                 
                 23246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100110; B = 8'b00000001; // Expected: {'P': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100110; B = 8'b00000001; | Outputs: P=%b | Expected: P=%d",
                 498,
                 
                 P
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010000; B = 8'b01111111; // Expected: {'P': 2032}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010000; B = 8'b01111111; | Outputs: P=%b | Expected: P=%d",
                 499,
                 
                 P
                 , 
                 
                 2032
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010101; B = 8'b11101010; // Expected: {'P': 4914}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010101; B = 8'b11101010; | Outputs: P=%b | Expected: P=%d",
                 500,
                 
                 P
                 , 
                 
                 4914
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111000; B = 8'b10100010; // Expected: {'P': 9072}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111000; B = 8'b10100010; | Outputs: P=%b | Expected: P=%d",
                 501,
                 
                 P
                 , 
                 
                 9072
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010011; B = 8'b11010001; // Expected: {'P': 17347}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010011; B = 8'b11010001; | Outputs: P=%b | Expected: P=%d",
                 502,
                 
                 P
                 , 
                 
                 17347
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010011; B = 8'b01011100; // Expected: {'P': 1748}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010011; B = 8'b01011100; | Outputs: P=%b | Expected: P=%d",
                 503,
                 
                 P
                 , 
                 
                 1748
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110111; B = 8'b11110001; // Expected: {'P': 28679}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110111; B = 8'b11110001; | Outputs: P=%b | Expected: P=%d",
                 504,
                 
                 P
                 , 
                 
                 28679
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100101; B = 8'b11101011; // Expected: {'P': 23735}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100101; B = 8'b11101011; | Outputs: P=%b | Expected: P=%d",
                 505,
                 
                 P
                 , 
                 
                 23735
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111001; B = 8'b11001011; // Expected: {'P': 24563}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111001; B = 8'b11001011; | Outputs: P=%b | Expected: P=%d",
                 506,
                 
                 P
                 , 
                 
                 24563
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100010; B = 8'b00100101; // Expected: {'P': 5994}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100010; B = 8'b00100101; | Outputs: P=%b | Expected: P=%d",
                 507,
                 
                 P
                 , 
                 
                 5994
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100011; B = 8'b01111110; // Expected: {'P': 4410}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100011; B = 8'b01111110; | Outputs: P=%b | Expected: P=%d",
                 508,
                 
                 P
                 , 
                 
                 4410
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111101; B = 8'b00110111; // Expected: {'P': 3355}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111101; B = 8'b00110111; | Outputs: P=%b | Expected: P=%d",
                 509,
                 
                 P
                 , 
                 
                 3355
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011011; B = 8'b11000111; // Expected: {'P': 30845}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011011; B = 8'b11000111; | Outputs: P=%b | Expected: P=%d",
                 510,
                 
                 P
                 , 
                 
                 30845
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001011; B = 8'b00111100; // Expected: {'P': 8340}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001011; B = 8'b00111100; | Outputs: P=%b | Expected: P=%d",
                 511,
                 
                 P
                 , 
                 
                 8340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110100; B = 8'b10001011; // Expected: {'P': 33916}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110100; B = 8'b10001011; | Outputs: P=%b | Expected: P=%d",
                 512,
                 
                 P
                 , 
                 
                 33916
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101010; B = 8'b10111111; // Expected: {'P': 8022}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101010; B = 8'b10111111; | Outputs: P=%b | Expected: P=%d",
                 513,
                 
                 P
                 , 
                 
                 8022
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100000; B = 8'b10101000; // Expected: {'P': 16128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100000; B = 8'b10101000; | Outputs: P=%b | Expected: P=%d",
                 514,
                 
                 P
                 , 
                 
                 16128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000101; B = 8'b10010101; // Expected: {'P': 745}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000101; B = 8'b10010101; | Outputs: P=%b | Expected: P=%d",
                 515,
                 
                 P
                 , 
                 
                 745
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100010; B = 8'b01100100; // Expected: {'P': 16200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100010; B = 8'b01100100; | Outputs: P=%b | Expected: P=%d",
                 516,
                 
                 P
                 , 
                 
                 16200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000100; B = 8'b10000011; // Expected: {'P': 17292}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000100; B = 8'b10000011; | Outputs: P=%b | Expected: P=%d",
                 517,
                 
                 P
                 , 
                 
                 17292
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101100; B = 8'b01110000; // Expected: {'P': 19264}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101100; B = 8'b01110000; | Outputs: P=%b | Expected: P=%d",
                 518,
                 
                 P
                 , 
                 
                 19264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111101; B = 8'b10111010; // Expected: {'P': 23250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111101; B = 8'b10111010; | Outputs: P=%b | Expected: P=%d",
                 519,
                 
                 P
                 , 
                 
                 23250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011010; B = 8'b00100011; // Expected: {'P': 3150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011010; B = 8'b00100011; | Outputs: P=%b | Expected: P=%d",
                 520,
                 
                 P
                 , 
                 
                 3150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111101; B = 8'b10000000; // Expected: {'P': 16000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111101; B = 8'b10000000; | Outputs: P=%b | Expected: P=%d",
                 521,
                 
                 P
                 , 
                 
                 16000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101010; B = 8'b01001100; // Expected: {'P': 12920}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101010; B = 8'b01001100; | Outputs: P=%b | Expected: P=%d",
                 522,
                 
                 P
                 , 
                 
                 12920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010000; B = 8'b00001100; // Expected: {'P': 960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010000; B = 8'b00001100; | Outputs: P=%b | Expected: P=%d",
                 523,
                 
                 P
                 , 
                 
                 960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011110; B = 8'b10011010; // Expected: {'P': 34188}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011110; B = 8'b10011010; | Outputs: P=%b | Expected: P=%d",
                 524,
                 
                 P
                 , 
                 
                 34188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110011; B = 8'b10110001; // Expected: {'P': 43011}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110011; B = 8'b10110001; | Outputs: P=%b | Expected: P=%d",
                 525,
                 
                 P
                 , 
                 
                 43011
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000011; B = 8'b10111011; // Expected: {'P': 12529}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000011; B = 8'b10111011; | Outputs: P=%b | Expected: P=%d",
                 526,
                 
                 P
                 , 
                 
                 12529
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001000; B = 8'b11010101; // Expected: {'P': 42600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001000; B = 8'b11010101; | Outputs: P=%b | Expected: P=%d",
                 527,
                 
                 P
                 , 
                 
                 42600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011101; B = 8'b10010101; // Expected: {'P': 32929}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011101; B = 8'b10010101; | Outputs: P=%b | Expected: P=%d",
                 528,
                 
                 P
                 , 
                 
                 32929
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001111; B = 8'b11101001; // Expected: {'P': 48231}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001111; B = 8'b11101001; | Outputs: P=%b | Expected: P=%d",
                 529,
                 
                 P
                 , 
                 
                 48231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000100; B = 8'b01101001; // Expected: {'P': 13860}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000100; B = 8'b01101001; | Outputs: P=%b | Expected: P=%d",
                 530,
                 
                 P
                 , 
                 
                 13860
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001000; B = 8'b11000001; // Expected: {'P': 26248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001000; B = 8'b11000001; | Outputs: P=%b | Expected: P=%d",
                 531,
                 
                 P
                 , 
                 
                 26248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000001; B = 8'b10110111; // Expected: {'P': 35319}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000001; B = 8'b10110111; | Outputs: P=%b | Expected: P=%d",
                 532,
                 
                 P
                 , 
                 
                 35319
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010101; B = 8'b00001111; // Expected: {'P': 2235}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010101; B = 8'b00001111; | Outputs: P=%b | Expected: P=%d",
                 533,
                 
                 P
                 , 
                 
                 2235
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010001; B = 8'b10110010; // Expected: {'P': 14418}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010001; B = 8'b10110010; | Outputs: P=%b | Expected: P=%d",
                 534,
                 
                 P
                 , 
                 
                 14418
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110100; B = 8'b00010010; // Expected: {'P': 4392}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110100; B = 8'b00010010; | Outputs: P=%b | Expected: P=%d",
                 535,
                 
                 P
                 , 
                 
                 4392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011001; B = 8'b01001111; // Expected: {'P': 1975}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011001; B = 8'b01001111; | Outputs: P=%b | Expected: P=%d",
                 536,
                 
                 P
                 , 
                 
                 1975
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100011; B = 8'b00010000; // Expected: {'P': 560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100011; B = 8'b00010000; | Outputs: P=%b | Expected: P=%d",
                 537,
                 
                 P
                 , 
                 
                 560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010001; B = 8'b10111001; // Expected: {'P': 14985}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010001; B = 8'b10111001; | Outputs: P=%b | Expected: P=%d",
                 538,
                 
                 P
                 , 
                 
                 14985
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001000; B = 8'b11111111; // Expected: {'P': 51000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001000; B = 8'b11111111; | Outputs: P=%b | Expected: P=%d",
                 539,
                 
                 P
                 , 
                 
                 51000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000011; B = 8'b10001111; // Expected: {'P': 18733}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000011; B = 8'b10001111; | Outputs: P=%b | Expected: P=%d",
                 540,
                 
                 P
                 , 
                 
                 18733
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110100; B = 8'b11111011; // Expected: {'P': 29116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110100; B = 8'b11111011; | Outputs: P=%b | Expected: P=%d",
                 541,
                 
                 P
                 , 
                 
                 29116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011000; B = 8'b00011110; // Expected: {'P': 4560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011000; B = 8'b00011110; | Outputs: P=%b | Expected: P=%d",
                 542,
                 
                 P
                 , 
                 
                 4560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011000; B = 8'b11011011; // Expected: {'P': 47304}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011000; B = 8'b11011011; | Outputs: P=%b | Expected: P=%d",
                 543,
                 
                 P
                 , 
                 
                 47304
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111110; B = 8'b00011110; // Expected: {'P': 5700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111110; B = 8'b00011110; | Outputs: P=%b | Expected: P=%d",
                 544,
                 
                 P
                 , 
                 
                 5700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100010; B = 8'b10010010; // Expected: {'P': 14308}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100010; B = 8'b10010010; | Outputs: P=%b | Expected: P=%d",
                 545,
                 
                 P
                 , 
                 
                 14308
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000011; B = 8'b00110111; // Expected: {'P': 165}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000011; B = 8'b00110111; | Outputs: P=%b | Expected: P=%d",
                 546,
                 
                 P
                 , 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111111; B = 8'b00011110; // Expected: {'P': 7650}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111111; B = 8'b00011110; | Outputs: P=%b | Expected: P=%d",
                 547,
                 
                 P
                 , 
                 
                 7650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110100; B = 8'b11011011; // Expected: {'P': 53436}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110100; B = 8'b11011011; | Outputs: P=%b | Expected: P=%d",
                 548,
                 
                 P
                 , 
                 
                 53436
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010000; B = 8'b00000111; // Expected: {'P': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010000; B = 8'b00000111; | Outputs: P=%b | Expected: P=%d",
                 549,
                 
                 P
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110110; B = 8'b10011111; // Expected: {'P': 8586}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110110; B = 8'b10011111; | Outputs: P=%b | Expected: P=%d",
                 550,
                 
                 P
                 , 
                 
                 8586
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100010; B = 8'b00101001; // Expected: {'P': 1394}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100010; B = 8'b00101001; | Outputs: P=%b | Expected: P=%d",
                 551,
                 
                 P
                 , 
                 
                 1394
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101011; B = 8'b10111111; // Expected: {'P': 32661}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101011; B = 8'b10111111; | Outputs: P=%b | Expected: P=%d",
                 552,
                 
                 P
                 , 
                 
                 32661
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110111; B = 8'b01101111; // Expected: {'P': 13209}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110111; B = 8'b01101111; | Outputs: P=%b | Expected: P=%d",
                 553,
                 
                 P
                 , 
                 
                 13209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100001; B = 8'b11100010; // Expected: {'P': 36386}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100001; B = 8'b11100010; | Outputs: P=%b | Expected: P=%d",
                 554,
                 
                 P
                 , 
                 
                 36386
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111011; B = 8'b10110110; // Expected: {'P': 45682}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111011; B = 8'b10110110; | Outputs: P=%b | Expected: P=%d",
                 555,
                 
                 P
                 , 
                 
                 45682
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100000; B = 8'b00001110; // Expected: {'P': 2240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100000; B = 8'b00001110; | Outputs: P=%b | Expected: P=%d",
                 556,
                 
                 P
                 , 
                 
                 2240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000110; B = 8'b10100001; // Expected: {'P': 31878}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000110; B = 8'b10100001; | Outputs: P=%b | Expected: P=%d",
                 557,
                 
                 P
                 , 
                 
                 31878
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001010; B = 8'b01011001; // Expected: {'P': 12282}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001010; B = 8'b01011001; | Outputs: P=%b | Expected: P=%d",
                 558,
                 
                 P
                 , 
                 
                 12282
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001110; B = 8'b01111010; // Expected: {'P': 17324}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001110; B = 8'b01111010; | Outputs: P=%b | Expected: P=%d",
                 559,
                 
                 P
                 , 
                 
                 17324
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110000; B = 8'b00001111; // Expected: {'P': 1680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110000; B = 8'b00001111; | Outputs: P=%b | Expected: P=%d",
                 560,
                 
                 P
                 , 
                 
                 1680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110100; B = 8'b00000010; // Expected: {'P': 360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110100; B = 8'b00000010; | Outputs: P=%b | Expected: P=%d",
                 561,
                 
                 P
                 , 
                 
                 360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011101; B = 8'b10000001; // Expected: {'P': 11997}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011101; B = 8'b10000001; | Outputs: P=%b | Expected: P=%d",
                 562,
                 
                 P
                 , 
                 
                 11997
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000100; B = 8'b01111011; // Expected: {'P': 8364}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000100; B = 8'b01111011; | Outputs: P=%b | Expected: P=%d",
                 563,
                 
                 P
                 , 
                 
                 8364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101001; B = 8'b11100111; // Expected: {'P': 39039}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101001; B = 8'b11100111; | Outputs: P=%b | Expected: P=%d",
                 564,
                 
                 P
                 , 
                 
                 39039
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110110; B = 8'b01010110; // Expected: {'P': 10148}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110110; B = 8'b01010110; | Outputs: P=%b | Expected: P=%d",
                 565,
                 
                 P
                 , 
                 
                 10148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100000; B = 8'b11000100; // Expected: {'P': 6272}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100000; B = 8'b11000100; | Outputs: P=%b | Expected: P=%d",
                 566,
                 
                 P
                 , 
                 
                 6272
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000000; B = 8'b01010010; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000000; B = 8'b01010010; | Outputs: P=%b | Expected: P=%d",
                 567,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000110; B = 8'b11011111; // Expected: {'P': 44154}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000110; B = 8'b11011111; | Outputs: P=%b | Expected: P=%d",
                 568,
                 
                 P
                 , 
                 
                 44154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101110; B = 8'b11001110; // Expected: {'P': 49028}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101110; B = 8'b11001110; | Outputs: P=%b | Expected: P=%d",
                 569,
                 
                 P
                 , 
                 
                 49028
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101110; B = 8'b01011000; // Expected: {'P': 9680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101110; B = 8'b01011000; | Outputs: P=%b | Expected: P=%d",
                 570,
                 
                 P
                 , 
                 
                 9680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101011; B = 8'b11000101; // Expected: {'P': 33687}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101011; B = 8'b11000101; | Outputs: P=%b | Expected: P=%d",
                 571,
                 
                 P
                 , 
                 
                 33687
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001011; B = 8'b00011100; // Expected: {'P': 308}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001011; B = 8'b00011100; | Outputs: P=%b | Expected: P=%d",
                 572,
                 
                 P
                 , 
                 
                 308
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101000; B = 8'b11000110; // Expected: {'P': 7920}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101000; B = 8'b11000110; | Outputs: P=%b | Expected: P=%d",
                 573,
                 
                 P
                 , 
                 
                 7920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010000; B = 8'b10110011; // Expected: {'P': 25776}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010000; B = 8'b10110011; | Outputs: P=%b | Expected: P=%d",
                 574,
                 
                 P
                 , 
                 
                 25776
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000010; B = 8'b11000011; // Expected: {'P': 390}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000010; B = 8'b11000011; | Outputs: P=%b | Expected: P=%d",
                 575,
                 
                 P
                 , 
                 
                 390
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010001; B = 8'b10101111; // Expected: {'P': 14175}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010001; B = 8'b10101111; | Outputs: P=%b | Expected: P=%d",
                 576,
                 
                 P
                 , 
                 
                 14175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100100; B = 8'b00010100; // Expected: {'P': 2000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100100; B = 8'b00010100; | Outputs: P=%b | Expected: P=%d",
                 577,
                 
                 P
                 , 
                 
                 2000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110111; B = 8'b01100111; // Expected: {'P': 18849}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110111; B = 8'b01100111; | Outputs: P=%b | Expected: P=%d",
                 578,
                 
                 P
                 , 
                 
                 18849
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101100; B = 8'b11010000; // Expected: {'P': 35776}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101100; B = 8'b11010000; | Outputs: P=%b | Expected: P=%d",
                 579,
                 
                 P
                 , 
                 
                 35776
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010101; B = 8'b11010010; // Expected: {'P': 4410}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010101; B = 8'b11010010; | Outputs: P=%b | Expected: P=%d",
                 580,
                 
                 P
                 , 
                 
                 4410
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011011; B = 8'b00000110; // Expected: {'P': 1314}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011011; B = 8'b00000110; | Outputs: P=%b | Expected: P=%d",
                 581,
                 
                 P
                 , 
                 
                 1314
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100100; B = 8'b01100000; // Expected: {'P': 21888}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100100; B = 8'b01100000; | Outputs: P=%b | Expected: P=%d",
                 582,
                 
                 P
                 , 
                 
                 21888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000000; B = 8'b10100101; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000000; B = 8'b10100101; | Outputs: P=%b | Expected: P=%d",
                 583,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010010; B = 8'b00100111; // Expected: {'P': 3198}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010010; B = 8'b00100111; | Outputs: P=%b | Expected: P=%d",
                 584,
                 
                 P
                 , 
                 
                 3198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101001; B = 8'b01100010; // Expected: {'P': 22834}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101001; B = 8'b01100010; | Outputs: P=%b | Expected: P=%d",
                 585,
                 
                 P
                 , 
                 
                 22834
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110110; B = 8'b11010011; // Expected: {'P': 51906}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110110; B = 8'b11010011; | Outputs: P=%b | Expected: P=%d",
                 586,
                 
                 P
                 , 
                 
                 51906
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000010; B = 8'b00110000; // Expected: {'P': 6240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000010; B = 8'b00110000; | Outputs: P=%b | Expected: P=%d",
                 587,
                 
                 P
                 , 
                 
                 6240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000000; B = 8'b00110101; // Expected: {'P': 3392}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000000; B = 8'b00110101; | Outputs: P=%b | Expected: P=%d",
                 588,
                 
                 P
                 , 
                 
                 3392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100100; B = 8'b10111110; // Expected: {'P': 6840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100100; B = 8'b10111110; | Outputs: P=%b | Expected: P=%d",
                 589,
                 
                 P
                 , 
                 
                 6840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110110; B = 8'b01001001; // Expected: {'P': 13286}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110110; B = 8'b01001001; | Outputs: P=%b | Expected: P=%d",
                 590,
                 
                 P
                 , 
                 
                 13286
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010010; B = 8'b01111001; // Expected: {'P': 2178}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010010; B = 8'b01111001; | Outputs: P=%b | Expected: P=%d",
                 591,
                 
                 P
                 , 
                 
                 2178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101011; B = 8'b01010010; // Expected: {'P': 8774}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101011; B = 8'b01010010; | Outputs: P=%b | Expected: P=%d",
                 592,
                 
                 P
                 , 
                 
                 8774
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100110; B = 8'b11100000; // Expected: {'P': 37184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100110; B = 8'b11100000; | Outputs: P=%b | Expected: P=%d",
                 593,
                 
                 P
                 , 
                 
                 37184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000101; B = 8'b10001001; // Expected: {'P': 9453}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000101; B = 8'b10001001; | Outputs: P=%b | Expected: P=%d",
                 594,
                 
                 P
                 , 
                 
                 9453
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101110; B = 8'b11011011; // Expected: {'P': 24090}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101110; B = 8'b11011011; | Outputs: P=%b | Expected: P=%d",
                 595,
                 
                 P
                 , 
                 
                 24090
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001000; B = 8'b10100111; // Expected: {'P': 1336}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001000; B = 8'b10100111; | Outputs: P=%b | Expected: P=%d",
                 596,
                 
                 P
                 , 
                 
                 1336
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100001; B = 8'b00000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100001; B = 8'b00000000; | Outputs: P=%b | Expected: P=%d",
                 597,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101011; B = 8'b10001010; // Expected: {'P': 14766}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101011; B = 8'b10001010; | Outputs: P=%b | Expected: P=%d",
                 598,
                 
                 P
                 , 
                 
                 14766
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000010; B = 8'b00110001; // Expected: {'P': 9506}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000010; B = 8'b00110001; | Outputs: P=%b | Expected: P=%d",
                 599,
                 
                 P
                 , 
                 
                 9506
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110110; B = 8'b00110111; // Expected: {'P': 10010}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110110; B = 8'b00110111; | Outputs: P=%b | Expected: P=%d",
                 600,
                 
                 P
                 , 
                 
                 10010
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110101; B = 8'b11101000; // Expected: {'P': 41992}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110101; B = 8'b11101000; | Outputs: P=%b | Expected: P=%d",
                 601,
                 
                 P
                 , 
                 
                 41992
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101100; B = 8'b11100100; // Expected: {'P': 10032}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101100; B = 8'b11100100; | Outputs: P=%b | Expected: P=%d",
                 602,
                 
                 P
                 , 
                 
                 10032
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001101; B = 8'b01001001; // Expected: {'P': 5621}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001101; B = 8'b01001001; | Outputs: P=%b | Expected: P=%d",
                 603,
                 
                 P
                 , 
                 
                 5621
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010100; B = 8'b11011111; // Expected: {'P': 33004}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010100; B = 8'b11011111; | Outputs: P=%b | Expected: P=%d",
                 604,
                 
                 P
                 , 
                 
                 33004
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001101; B = 8'b01000010; // Expected: {'P': 858}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001101; B = 8'b01000010; | Outputs: P=%b | Expected: P=%d",
                 605,
                 
                 P
                 , 
                 
                 858
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010101; B = 8'b11101100; // Expected: {'P': 4956}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010101; B = 8'b11101100; | Outputs: P=%b | Expected: P=%d",
                 606,
                 
                 P
                 , 
                 
                 4956
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111111; B = 8'b11111011; // Expected: {'P': 47941}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111111; B = 8'b11111011; | Outputs: P=%b | Expected: P=%d",
                 607,
                 
                 P
                 , 
                 
                 47941
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001110; B = 8'b10111100; // Expected: {'P': 26696}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001110; B = 8'b10111100; | Outputs: P=%b | Expected: P=%d",
                 608,
                 
                 P
                 , 
                 
                 26696
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001110; B = 8'b01001011; // Expected: {'P': 1050}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001110; B = 8'b01001011; | Outputs: P=%b | Expected: P=%d",
                 609,
                 
                 P
                 , 
                 
                 1050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000010; B = 8'b00010111; // Expected: {'P': 4462}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000010; B = 8'b00010111; | Outputs: P=%b | Expected: P=%d",
                 610,
                 
                 P
                 , 
                 
                 4462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101100; B = 8'b00111010; // Expected: {'P': 13688}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101100; B = 8'b00111010; | Outputs: P=%b | Expected: P=%d",
                 611,
                 
                 P
                 , 
                 
                 13688
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000100; B = 8'b10100001; // Expected: {'P': 31556}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000100; B = 8'b10100001; | Outputs: P=%b | Expected: P=%d",
                 612,
                 
                 P
                 , 
                 
                 31556
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000111; B = 8'b11110000; // Expected: {'P': 47760}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000111; B = 8'b11110000; | Outputs: P=%b | Expected: P=%d",
                 613,
                 
                 P
                 , 
                 
                 47760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001111; B = 8'b10011010; // Expected: {'P': 12166}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001111; B = 8'b10011010; | Outputs: P=%b | Expected: P=%d",
                 614,
                 
                 P
                 , 
                 
                 12166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010110; B = 8'b00101110; // Expected: {'P': 3956}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010110; B = 8'b00101110; | Outputs: P=%b | Expected: P=%d",
                 615,
                 
                 P
                 , 
                 
                 3956
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001010; B = 8'b00011111; // Expected: {'P': 2294}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001010; B = 8'b00011111; | Outputs: P=%b | Expected: P=%d",
                 616,
                 
                 P
                 , 
                 
                 2294
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110100; B = 8'b01010000; // Expected: {'P': 9280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110100; B = 8'b01010000; | Outputs: P=%b | Expected: P=%d",
                 617,
                 
                 P
                 , 
                 
                 9280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100011; B = 8'b00001100; // Expected: {'P': 1188}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100011; B = 8'b00001100; | Outputs: P=%b | Expected: P=%d",
                 618,
                 
                 P
                 , 
                 
                 1188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110011; B = 8'b01001001; // Expected: {'P': 3723}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110011; B = 8'b01001001; | Outputs: P=%b | Expected: P=%d",
                 619,
                 
                 P
                 , 
                 
                 3723
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110010; B = 8'b00010010; // Expected: {'P': 2052}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110010; B = 8'b00010010; | Outputs: P=%b | Expected: P=%d",
                 620,
                 
                 P
                 , 
                 
                 2052
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011001; B = 8'b00011100; // Expected: {'P': 2492}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011001; B = 8'b00011100; | Outputs: P=%b | Expected: P=%d",
                 621,
                 
                 P
                 , 
                 
                 2492
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000000; B = 8'b00011001; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000000; B = 8'b00011001; | Outputs: P=%b | Expected: P=%d",
                 622,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011001; B = 8'b00101101; // Expected: {'P': 6885}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011001; B = 8'b00101101; | Outputs: P=%b | Expected: P=%d",
                 623,
                 
                 P
                 , 
                 
                 6885
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000100; B = 8'b01010111; // Expected: {'P': 5916}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000100; B = 8'b01010111; | Outputs: P=%b | Expected: P=%d",
                 624,
                 
                 P
                 , 
                 
                 5916
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011101; B = 8'b10011000; // Expected: {'P': 4408}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011101; B = 8'b10011000; | Outputs: P=%b | Expected: P=%d",
                 625,
                 
                 P
                 , 
                 
                 4408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100101; B = 8'b01110110; // Expected: {'P': 19470}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100101; B = 8'b01110110; | Outputs: P=%b | Expected: P=%d",
                 626,
                 
                 P
                 , 
                 
                 19470
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000011; B = 8'b00011110; // Expected: {'P': 5850}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000011; B = 8'b00011110; | Outputs: P=%b | Expected: P=%d",
                 627,
                 
                 P
                 , 
                 
                 5850
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111010; B = 8'b11101001; // Expected: {'P': 58250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111010; B = 8'b11101001; | Outputs: P=%b | Expected: P=%d",
                 628,
                 
                 P
                 , 
                 
                 58250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111010; B = 8'b01000000; // Expected: {'P': 3712}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111010; B = 8'b01000000; | Outputs: P=%b | Expected: P=%d",
                 629,
                 
                 P
                 , 
                 
                 3712
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100110; B = 8'b10010100; // Expected: {'P': 15096}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100110; B = 8'b10010100; | Outputs: P=%b | Expected: P=%d",
                 630,
                 
                 P
                 , 
                 
                 15096
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001001; B = 8'b00100100; // Expected: {'P': 4932}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001001; B = 8'b00100100; | Outputs: P=%b | Expected: P=%d",
                 631,
                 
                 P
                 , 
                 
                 4932
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100100; B = 8'b00100110; // Expected: {'P': 8664}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100100; B = 8'b00100110; | Outputs: P=%b | Expected: P=%d",
                 632,
                 
                 P
                 , 
                 
                 8664
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101111; B = 8'b11000111; // Expected: {'P': 22089}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101111; B = 8'b11000111; | Outputs: P=%b | Expected: P=%d",
                 633,
                 
                 P
                 , 
                 
                 22089
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100100; B = 8'b00111111; // Expected: {'P': 6300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100100; B = 8'b00111111; | Outputs: P=%b | Expected: P=%d",
                 634,
                 
                 P
                 , 
                 
                 6300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100010; B = 8'b00010110; // Expected: {'P': 748}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100010; B = 8'b00010110; | Outputs: P=%b | Expected: P=%d",
                 635,
                 
                 P
                 , 
                 
                 748
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111011; B = 8'b11000010; // Expected: {'P': 11446}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111011; B = 8'b11000010; | Outputs: P=%b | Expected: P=%d",
                 636,
                 
                 P
                 , 
                 
                 11446
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000000; B = 8'b00011111; // Expected: {'P': 3968}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000000; B = 8'b00011111; | Outputs: P=%b | Expected: P=%d",
                 637,
                 
                 P
                 , 
                 
                 3968
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001001; B = 8'b11010111; // Expected: {'P': 1935}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001001; B = 8'b11010111; | Outputs: P=%b | Expected: P=%d",
                 638,
                 
                 P
                 , 
                 
                 1935
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011100; B = 8'b11000110; // Expected: {'P': 43560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011100; B = 8'b11000110; | Outputs: P=%b | Expected: P=%d",
                 639,
                 
                 P
                 , 
                 
                 43560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110011; B = 8'b00001010; // Expected: {'P': 1150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110011; B = 8'b00001010; | Outputs: P=%b | Expected: P=%d",
                 640,
                 
                 P
                 , 
                 
                 1150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100000; B = 8'b01101010; // Expected: {'P': 10176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100000; B = 8'b01101010; | Outputs: P=%b | Expected: P=%d",
                 641,
                 
                 P
                 , 
                 
                 10176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000000; B = 8'b01100101; // Expected: {'P': 12928}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000000; B = 8'b01100101; | Outputs: P=%b | Expected: P=%d",
                 642,
                 
                 P
                 , 
                 
                 12928
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000101; B = 8'b11011000; // Expected: {'P': 14904}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000101; B = 8'b11011000; | Outputs: P=%b | Expected: P=%d",
                 643,
                 
                 P
                 , 
                 
                 14904
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100010; B = 8'b01101010; // Expected: {'P': 17172}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100010; B = 8'b01101010; | Outputs: P=%b | Expected: P=%d",
                 644,
                 
                 P
                 , 
                 
                 17172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111101; B = 8'b01000000; // Expected: {'P': 8000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111101; B = 8'b01000000; | Outputs: P=%b | Expected: P=%d",
                 645,
                 
                 P
                 , 
                 
                 8000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100101; B = 8'b10001111; // Expected: {'P': 5291}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100101; B = 8'b10001111; | Outputs: P=%b | Expected: P=%d",
                 646,
                 
                 P
                 , 
                 
                 5291
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000010; B = 8'b01100011; // Expected: {'P': 198}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000010; B = 8'b01100011; | Outputs: P=%b | Expected: P=%d",
                 647,
                 
                 P
                 , 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100111; B = 8'b01110100; // Expected: {'P': 4524}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100111; B = 8'b01110100; | Outputs: P=%b | Expected: P=%d",
                 648,
                 
                 P
                 , 
                 
                 4524
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111011; B = 8'b01101011; // Expected: {'P': 20009}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111011; B = 8'b01101011; | Outputs: P=%b | Expected: P=%d",
                 649,
                 
                 P
                 , 
                 
                 20009
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010000; B = 8'b11111110; // Expected: {'P': 52832}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010000; B = 8'b11111110; | Outputs: P=%b | Expected: P=%d",
                 650,
                 
                 P
                 , 
                 
                 52832
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010100; B = 8'b10000011; // Expected: {'P': 19388}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010100; B = 8'b10000011; | Outputs: P=%b | Expected: P=%d",
                 651,
                 
                 P
                 , 
                 
                 19388
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100110; B = 8'b11010111; // Expected: {'P': 21930}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100110; B = 8'b11010111; | Outputs: P=%b | Expected: P=%d",
                 652,
                 
                 P
                 , 
                 
                 21930
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100010; B = 8'b11101110; // Expected: {'P': 53788}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100010; B = 8'b11101110; | Outputs: P=%b | Expected: P=%d",
                 653,
                 
                 P
                 , 
                 
                 53788
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100010; B = 8'b01010111; // Expected: {'P': 2958}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100010; B = 8'b01010111; | Outputs: P=%b | Expected: P=%d",
                 654,
                 
                 P
                 , 
                 
                 2958
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100110; B = 8'b00110000; // Expected: {'P': 1824}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100110; B = 8'b00110000; | Outputs: P=%b | Expected: P=%d",
                 655,
                 
                 P
                 , 
                 
                 1824
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111111; B = 8'b10101110; // Expected: {'P': 33234}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111111; B = 8'b10101110; | Outputs: P=%b | Expected: P=%d",
                 656,
                 
                 P
                 , 
                 
                 33234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110000; B = 8'b11010101; // Expected: {'P': 37488}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110000; B = 8'b11010101; | Outputs: P=%b | Expected: P=%d",
                 657,
                 
                 P
                 , 
                 
                 37488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101010; B = 8'b00011010; // Expected: {'P': 2756}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101010; B = 8'b00011010; | Outputs: P=%b | Expected: P=%d",
                 658,
                 
                 P
                 , 
                 
                 2756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100001; B = 8'b00110001; // Expected: {'P': 7889}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100001; B = 8'b00110001; | Outputs: P=%b | Expected: P=%d",
                 659,
                 
                 P
                 , 
                 
                 7889
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111011; B = 8'b10001100; // Expected: {'P': 8260}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111011; B = 8'b10001100; | Outputs: P=%b | Expected: P=%d",
                 660,
                 
                 P
                 , 
                 
                 8260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110101; B = 8'b10011000; // Expected: {'P': 17784}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110101; B = 8'b10011000; | Outputs: P=%b | Expected: P=%d",
                 661,
                 
                 P
                 , 
                 
                 17784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111010; B = 8'b11111011; // Expected: {'P': 30622}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111010; B = 8'b11111011; | Outputs: P=%b | Expected: P=%d",
                 662,
                 
                 P
                 , 
                 
                 30622
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110001; B = 8'b11101111; // Expected: {'P': 42303}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110001; B = 8'b11101111; | Outputs: P=%b | Expected: P=%d",
                 663,
                 
                 P
                 , 
                 
                 42303
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001100; B = 8'b01001110; // Expected: {'P': 10920}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001100; B = 8'b01001110; | Outputs: P=%b | Expected: P=%d",
                 664,
                 
                 P
                 , 
                 
                 10920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111010; B = 8'b11111101; // Expected: {'P': 14674}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111010; B = 8'b11111101; | Outputs: P=%b | Expected: P=%d",
                 665,
                 
                 P
                 , 
                 
                 14674
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110101; B = 8'b01101000; // Expected: {'P': 12168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110101; B = 8'b01101000; | Outputs: P=%b | Expected: P=%d",
                 666,
                 
                 P
                 , 
                 
                 12168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000101; B = 8'b00010111; // Expected: {'P': 115}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000101; B = 8'b00010111; | Outputs: P=%b | Expected: P=%d",
                 667,
                 
                 P
                 , 
                 
                 115
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100110; B = 8'b01000001; // Expected: {'P': 10790}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100110; B = 8'b01000001; | Outputs: P=%b | Expected: P=%d",
                 668,
                 
                 P
                 , 
                 
                 10790
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101011; B = 8'b00100111; // Expected: {'P': 1677}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101011; B = 8'b00100111; | Outputs: P=%b | Expected: P=%d",
                 669,
                 
                 P
                 , 
                 
                 1677
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000101; B = 8'b01000111; // Expected: {'P': 9443}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000101; B = 8'b01000111; | Outputs: P=%b | Expected: P=%d",
                 670,
                 
                 P
                 , 
                 
                 9443
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010111; B = 8'b01001000; // Expected: {'P': 10872}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010111; B = 8'b01001000; | Outputs: P=%b | Expected: P=%d",
                 671,
                 
                 P
                 , 
                 
                 10872
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010001; B = 8'b00010110; // Expected: {'P': 4598}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010001; B = 8'b00010110; | Outputs: P=%b | Expected: P=%d",
                 672,
                 
                 P
                 , 
                 
                 4598
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100111; B = 8'b00111100; // Expected: {'P': 2340}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100111; B = 8'b00111100; | Outputs: P=%b | Expected: P=%d",
                 673,
                 
                 P
                 , 
                 
                 2340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000101; B = 8'b10100111; // Expected: {'P': 835}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000101; B = 8'b10100111; | Outputs: P=%b | Expected: P=%d",
                 674,
                 
                 P
                 , 
                 
                 835
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011110; B = 8'b10010100; // Expected: {'P': 32856}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011110; B = 8'b10010100; | Outputs: P=%b | Expected: P=%d",
                 675,
                 
                 P
                 , 
                 
                 32856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110111; B = 8'b11001111; // Expected: {'P': 37881}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110111; B = 8'b11001111; | Outputs: P=%b | Expected: P=%d",
                 676,
                 
                 P
                 , 
                 
                 37881
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111100; B = 8'b01110110; // Expected: {'P': 22184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111100; B = 8'b01110110; | Outputs: P=%b | Expected: P=%d",
                 677,
                 
                 P
                 , 
                 
                 22184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101100; B = 8'b10100000; // Expected: {'P': 27520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101100; B = 8'b10100000; | Outputs: P=%b | Expected: P=%d",
                 678,
                 
                 P
                 , 
                 
                 27520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101111; B = 8'b01001000; // Expected: {'P': 7992}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101111; B = 8'b01001000; | Outputs: P=%b | Expected: P=%d",
                 679,
                 
                 P
                 , 
                 
                 7992
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100110; B = 8'b11110111; // Expected: {'P': 56810}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100110; B = 8'b11110111; | Outputs: P=%b | Expected: P=%d",
                 680,
                 
                 P
                 , 
                 
                 56810
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100010; B = 8'b00111100; // Expected: {'P': 2040}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100010; B = 8'b00111100; | Outputs: P=%b | Expected: P=%d",
                 681,
                 
                 P
                 , 
                 
                 2040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000010; B = 8'b01101000; // Expected: {'P': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000010; B = 8'b01101000; | Outputs: P=%b | Expected: P=%d",
                 682,
                 
                 P
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010100; B = 8'b00100100; // Expected: {'P': 3024}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010100; B = 8'b00100100; | Outputs: P=%b | Expected: P=%d",
                 683,
                 
                 P
                 , 
                 
                 3024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011001; B = 8'b01110100; // Expected: {'P': 25172}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011001; B = 8'b01110100; | Outputs: P=%b | Expected: P=%d",
                 684,
                 
                 P
                 , 
                 
                 25172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000110; B = 8'b11101100; // Expected: {'P': 46728}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000110; B = 8'b11101100; | Outputs: P=%b | Expected: P=%d",
                 685,
                 
                 P
                 , 
                 
                 46728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001111; B = 8'b10000110; // Expected: {'P': 2010}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001111; B = 8'b10000110; | Outputs: P=%b | Expected: P=%d",
                 686,
                 
                 P
                 , 
                 
                 2010
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011000; B = 8'b11010100; // Expected: {'P': 18656}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011000; B = 8'b11010100; | Outputs: P=%b | Expected: P=%d",
                 687,
                 
                 P
                 , 
                 
                 18656
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101000; B = 8'b11110000; // Expected: {'P': 55680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101000; B = 8'b11110000; | Outputs: P=%b | Expected: P=%d",
                 688,
                 
                 P
                 , 
                 
                 55680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110000; B = 8'b01101011; // Expected: {'P': 5136}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110000; B = 8'b01101011; | Outputs: P=%b | Expected: P=%d",
                 689,
                 
                 P
                 , 
                 
                 5136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100101; B = 8'b00000100; // Expected: {'P': 148}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100101; B = 8'b00000100; | Outputs: P=%b | Expected: P=%d",
                 690,
                 
                 P
                 , 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101000; B = 8'b00000101; // Expected: {'P': 520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101000; B = 8'b00000101; | Outputs: P=%b | Expected: P=%d",
                 691,
                 
                 P
                 , 
                 
                 520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011000; B = 8'b10101001; // Expected: {'P': 25688}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011000; B = 8'b10101001; | Outputs: P=%b | Expected: P=%d",
                 692,
                 
                 P
                 , 
                 
                 25688
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000101; B = 8'b11011110; // Expected: {'P': 43734}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000101; B = 8'b11011110; | Outputs: P=%b | Expected: P=%d",
                 693,
                 
                 P
                 , 
                 
                 43734
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000000; B = 8'b10110000; // Expected: {'P': 22528}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000000; B = 8'b10110000; | Outputs: P=%b | Expected: P=%d",
                 694,
                 
                 P
                 , 
                 
                 22528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001101; B = 8'b01000100; // Expected: {'P': 9588}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001101; B = 8'b01000100; | Outputs: P=%b | Expected: P=%d",
                 695,
                 
                 P
                 , 
                 
                 9588
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100001; B = 8'b01110001; // Expected: {'P': 18193}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100001; B = 8'b01110001; | Outputs: P=%b | Expected: P=%d",
                 696,
                 
                 P
                 , 
                 
                 18193
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111011; B = 8'b01000101; // Expected: {'P': 8487}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111011; B = 8'b01000101; | Outputs: P=%b | Expected: P=%d",
                 697,
                 
                 P
                 , 
                 
                 8487
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001110; B = 8'b01111010; // Expected: {'P': 1708}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001110; B = 8'b01111010; | Outputs: P=%b | Expected: P=%d",
                 698,
                 
                 P
                 , 
                 
                 1708
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110111; B = 8'b00100111; // Expected: {'P': 2145}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110111; B = 8'b00100111; | Outputs: P=%b | Expected: P=%d",
                 699,
                 
                 P
                 , 
                 
                 2145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101000; B = 8'b11011100; // Expected: {'P': 36960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101000; B = 8'b11011100; | Outputs: P=%b | Expected: P=%d",
                 700,
                 
                 P
                 , 
                 
                 36960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001000; B = 8'b00100010; // Expected: {'P': 272}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001000; B = 8'b00100010; | Outputs: P=%b | Expected: P=%d",
                 701,
                 
                 P
                 , 
                 
                 272
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110010; B = 8'b00011001; // Expected: {'P': 6050}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110010; B = 8'b00011001; | Outputs: P=%b | Expected: P=%d",
                 702,
                 
                 P
                 , 
                 
                 6050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001010; B = 8'b01100101; // Expected: {'P': 13938}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001010; B = 8'b01100101; | Outputs: P=%b | Expected: P=%d",
                 703,
                 
                 P
                 , 
                 
                 13938
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001100; B = 8'b00101001; // Expected: {'P': 8364}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001100; B = 8'b00101001; | Outputs: P=%b | Expected: P=%d",
                 704,
                 
                 P
                 , 
                 
                 8364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110101; B = 8'b00010111; // Expected: {'P': 4163}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110101; B = 8'b00010111; | Outputs: P=%b | Expected: P=%d",
                 705,
                 
                 P
                 , 
                 
                 4163
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001000; B = 8'b11010111; // Expected: {'P': 29240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001000; B = 8'b11010111; | Outputs: P=%b | Expected: P=%d",
                 706,
                 
                 P
                 , 
                 
                 29240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010110; B = 8'b00001110; // Expected: {'P': 1204}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010110; B = 8'b00001110; | Outputs: P=%b | Expected: P=%d",
                 707,
                 
                 P
                 , 
                 
                 1204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000011; B = 8'b11101001; // Expected: {'P': 699}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000011; B = 8'b11101001; | Outputs: P=%b | Expected: P=%d",
                 708,
                 
                 P
                 , 
                 
                 699
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100101; B = 8'b11101001; // Expected: {'P': 38445}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100101; B = 8'b11101001; | Outputs: P=%b | Expected: P=%d",
                 709,
                 
                 P
                 , 
                 
                 38445
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001110; B = 8'b01000101; // Expected: {'P': 966}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001110; B = 8'b01000101; | Outputs: P=%b | Expected: P=%d",
                 710,
                 
                 P
                 , 
                 
                 966
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101111; B = 8'b11111101; // Expected: {'P': 11891}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101111; B = 8'b11111101; | Outputs: P=%b | Expected: P=%d",
                 711,
                 
                 P
                 , 
                 
                 11891
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001111; B = 8'b11100001; // Expected: {'P': 46575}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001111; B = 8'b11100001; | Outputs: P=%b | Expected: P=%d",
                 712,
                 
                 P
                 , 
                 
                 46575
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110010; B = 8'b10101100; // Expected: {'P': 19608}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110010; B = 8'b10101100; | Outputs: P=%b | Expected: P=%d",
                 713,
                 
                 P
                 , 
                 
                 19608
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111001; B = 8'b00000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111001; B = 8'b00000000; | Outputs: P=%b | Expected: P=%d",
                 714,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010001; B = 8'b11101110; // Expected: {'P': 34510}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010001; B = 8'b11101110; | Outputs: P=%b | Expected: P=%d",
                 715,
                 
                 P
                 , 
                 
                 34510
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101000; B = 8'b01100101; // Expected: {'P': 16968}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101000; B = 8'b01100101; | Outputs: P=%b | Expected: P=%d",
                 716,
                 
                 P
                 , 
                 
                 16968
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101011; B = 8'b01101111; // Expected: {'P': 18981}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101011; B = 8'b01101111; | Outputs: P=%b | Expected: P=%d",
                 717,
                 
                 P
                 , 
                 
                 18981
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001001; B = 8'b11011110; // Expected: {'P': 1998}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001001; B = 8'b11011110; | Outputs: P=%b | Expected: P=%d",
                 718,
                 
                 P
                 , 
                 
                 1998
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011001; B = 8'b10001100; // Expected: {'P': 3500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011001; B = 8'b10001100; | Outputs: P=%b | Expected: P=%d",
                 719,
                 
                 P
                 , 
                 
                 3500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111010; B = 8'b10011000; // Expected: {'P': 8816}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111010; B = 8'b10011000; | Outputs: P=%b | Expected: P=%d",
                 720,
                 
                 P
                 , 
                 
                 8816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101011; B = 8'b11011001; // Expected: {'P': 9331}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101011; B = 8'b11011001; | Outputs: P=%b | Expected: P=%d",
                 721,
                 
                 P
                 , 
                 
                 9331
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001101; B = 8'b01110100; // Expected: {'P': 16356}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001101; B = 8'b01110100; | Outputs: P=%b | Expected: P=%d",
                 722,
                 
                 P
                 , 
                 
                 16356
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100000; B = 8'b11110110; // Expected: {'P': 55104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100000; B = 8'b11110110; | Outputs: P=%b | Expected: P=%d",
                 723,
                 
                 P
                 , 
                 
                 55104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101000; B = 8'b11001001; // Expected: {'P': 8040}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101000; B = 8'b11001001; | Outputs: P=%b | Expected: P=%d",
                 724,
                 
                 P
                 , 
                 
                 8040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110001; B = 8'b10001010; // Expected: {'P': 6762}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110001; B = 8'b10001010; | Outputs: P=%b | Expected: P=%d",
                 725,
                 
                 P
                 , 
                 
                 6762
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100010; B = 8'b00000111; // Expected: {'P': 686}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100010; B = 8'b00000111; | Outputs: P=%b | Expected: P=%d",
                 726,
                 
                 P
                 , 
                 
                 686
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100001; B = 8'b11010000; // Expected: {'P': 20176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100001; B = 8'b11010000; | Outputs: P=%b | Expected: P=%d",
                 727,
                 
                 P
                 , 
                 
                 20176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111111; B = 8'b01110100; // Expected: {'P': 29580}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111111; B = 8'b01110100; | Outputs: P=%b | Expected: P=%d",
                 728,
                 
                 P
                 , 
                 
                 29580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000110; B = 8'b10001110; // Expected: {'P': 852}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000110; B = 8'b10001110; | Outputs: P=%b | Expected: P=%d",
                 729,
                 
                 P
                 , 
                 
                 852
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110101; B = 8'b11101001; // Expected: {'P': 12349}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110101; B = 8'b11101001; | Outputs: P=%b | Expected: P=%d",
                 730,
                 
                 P
                 , 
                 
                 12349
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011100; B = 8'b00000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011100; B = 8'b00000000; | Outputs: P=%b | Expected: P=%d",
                 731,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101110; B = 8'b01000101; // Expected: {'P': 3174}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101110; B = 8'b01000101; | Outputs: P=%b | Expected: P=%d",
                 732,
                 
                 P
                 , 
                 
                 3174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101101; B = 8'b00000001; // Expected: {'P': 109}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101101; B = 8'b00000001; | Outputs: P=%b | Expected: P=%d",
                 733,
                 
                 P
                 , 
                 
                 109
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110100; B = 8'b10111001; // Expected: {'P': 21460}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110100; B = 8'b10111001; | Outputs: P=%b | Expected: P=%d",
                 734,
                 
                 P
                 , 
                 
                 21460
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101010; B = 8'b10011011; // Expected: {'P': 16430}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101010; B = 8'b10011011; | Outputs: P=%b | Expected: P=%d",
                 735,
                 
                 P
                 , 
                 
                 16430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100001; B = 8'b01111101; // Expected: {'P': 20125}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100001; B = 8'b01111101; | Outputs: P=%b | Expected: P=%d",
                 736,
                 
                 P
                 , 
                 
                 20125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001100; B = 8'b01101101; // Expected: {'P': 22236}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001100; B = 8'b01101101; | Outputs: P=%b | Expected: P=%d",
                 737,
                 
                 P
                 , 
                 
                 22236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100011; B = 8'b01001110; // Expected: {'P': 2730}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100011; B = 8'b01001110; | Outputs: P=%b | Expected: P=%d",
                 738,
                 
                 P
                 , 
                 
                 2730
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010110; B = 8'b01101100; // Expected: {'P': 23112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010110; B = 8'b01101100; | Outputs: P=%b | Expected: P=%d",
                 739,
                 
                 P
                 , 
                 
                 23112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101000; B = 8'b11100100; // Expected: {'P': 23712}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101000; B = 8'b11100100; | Outputs: P=%b | Expected: P=%d",
                 740,
                 
                 P
                 , 
                 
                 23712
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111011; B = 8'b11011001; // Expected: {'P': 26691}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111011; B = 8'b11011001; | Outputs: P=%b | Expected: P=%d",
                 741,
                 
                 P
                 , 
                 
                 26691
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011110; B = 8'b10000001; // Expected: {'P': 28638}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011110; B = 8'b10000001; | Outputs: P=%b | Expected: P=%d",
                 742,
                 
                 P
                 , 
                 
                 28638
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010001; B = 8'b11101010; // Expected: {'P': 48906}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010001; B = 8'b11101010; | Outputs: P=%b | Expected: P=%d",
                 743,
                 
                 P
                 , 
                 
                 48906
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100101; B = 8'b11000011; // Expected: {'P': 7215}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100101; B = 8'b11000011; | Outputs: P=%b | Expected: P=%d",
                 744,
                 
                 P
                 , 
                 
                 7215
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000001; B = 8'b10000111; // Expected: {'P': 135}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000001; B = 8'b10000111; | Outputs: P=%b | Expected: P=%d",
                 745,
                 
                 P
                 , 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101000; B = 8'b00100110; // Expected: {'P': 1520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101000; B = 8'b00100110; | Outputs: P=%b | Expected: P=%d",
                 746,
                 
                 P
                 , 
                 
                 1520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110000; B = 8'b10001010; // Expected: {'P': 33120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110000; B = 8'b10001010; | Outputs: P=%b | Expected: P=%d",
                 747,
                 
                 P
                 , 
                 
                 33120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001010; B = 8'b11101000; // Expected: {'P': 2320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001010; B = 8'b11101000; | Outputs: P=%b | Expected: P=%d",
                 748,
                 
                 P
                 , 
                 
                 2320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101110; B = 8'b11010110; // Expected: {'P': 50932}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101110; B = 8'b11010110; | Outputs: P=%b | Expected: P=%d",
                 749,
                 
                 P
                 , 
                 
                 50932
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010101; B = 8'b11010010; // Expected: {'P': 44730}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010101; B = 8'b11010010; | Outputs: P=%b | Expected: P=%d",
                 750,
                 
                 P
                 , 
                 
                 44730
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101110; B = 8'b00001000; // Expected: {'P': 1904}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101110; B = 8'b00001000; | Outputs: P=%b | Expected: P=%d",
                 751,
                 
                 P
                 , 
                 
                 1904
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010111; B = 8'b11001111; // Expected: {'P': 4761}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010111; B = 8'b11001111; | Outputs: P=%b | Expected: P=%d",
                 752,
                 
                 P
                 , 
                 
                 4761
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011111; B = 8'b10111110; // Expected: {'P': 18050}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011111; B = 8'b10111110; | Outputs: P=%b | Expected: P=%d",
                 753,
                 
                 P
                 , 
                 
                 18050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100110; B = 8'b01010101; // Expected: {'P': 3230}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100110; B = 8'b01010101; | Outputs: P=%b | Expected: P=%d",
                 754,
                 
                 P
                 , 
                 
                 3230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110010; B = 8'b11010101; // Expected: {'P': 10650}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110010; B = 8'b11010101; | Outputs: P=%b | Expected: P=%d",
                 755,
                 
                 P
                 , 
                 
                 10650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110101; B = 8'b10111001; // Expected: {'P': 9805}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110101; B = 8'b10111001; | Outputs: P=%b | Expected: P=%d",
                 756,
                 
                 P
                 , 
                 
                 9805
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100000; B = 8'b01011000; // Expected: {'P': 19712}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100000; B = 8'b01011000; | Outputs: P=%b | Expected: P=%d",
                 757,
                 
                 P
                 , 
                 
                 19712
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100011; B = 8'b11110001; // Expected: {'P': 54707}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100011; B = 8'b11110001; | Outputs: P=%b | Expected: P=%d",
                 758,
                 
                 P
                 , 
                 
                 54707
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010010; B = 8'b11000111; // Expected: {'P': 29054}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010010; B = 8'b11000111; | Outputs: P=%b | Expected: P=%d",
                 759,
                 
                 P
                 , 
                 
                 29054
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011110; B = 8'b10010011; // Expected: {'P': 32634}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011110; B = 8'b10010011; | Outputs: P=%b | Expected: P=%d",
                 760,
                 
                 P
                 , 
                 
                 32634
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110111; B = 8'b10111100; // Expected: {'P': 22372}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110111; B = 8'b10111100; | Outputs: P=%b | Expected: P=%d",
                 761,
                 
                 P
                 , 
                 
                 22372
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000010; B = 8'b10100011; // Expected: {'P': 21190}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000010; B = 8'b10100011; | Outputs: P=%b | Expected: P=%d",
                 762,
                 
                 P
                 , 
                 
                 21190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110100; B = 8'b01101100; // Expected: {'P': 26352}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110100; B = 8'b01101100; | Outputs: P=%b | Expected: P=%d",
                 763,
                 
                 P
                 , 
                 
                 26352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111110; B = 8'b10100001; // Expected: {'P': 9982}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111110; B = 8'b10100001; | Outputs: P=%b | Expected: P=%d",
                 764,
                 
                 P
                 , 
                 
                 9982
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001011; B = 8'b01010110; // Expected: {'P': 6450}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001011; B = 8'b01010110; | Outputs: P=%b | Expected: P=%d",
                 765,
                 
                 P
                 , 
                 
                 6450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000100; B = 8'b11000011; // Expected: {'P': 13260}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000100; B = 8'b11000011; | Outputs: P=%b | Expected: P=%d",
                 766,
                 
                 P
                 , 
                 
                 13260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101011; B = 8'b11111011; // Expected: {'P': 10793}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101011; B = 8'b11111011; | Outputs: P=%b | Expected: P=%d",
                 767,
                 
                 P
                 , 
                 
                 10793
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110111; B = 8'b00110011; // Expected: {'P': 12597}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110111; B = 8'b00110011; | Outputs: P=%b | Expected: P=%d",
                 768,
                 
                 P
                 , 
                 
                 12597
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011111; B = 8'b10000000; // Expected: {'P': 3968}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011111; B = 8'b10000000; | Outputs: P=%b | Expected: P=%d",
                 769,
                 
                 P
                 , 
                 
                 3968
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010101; B = 8'b10100000; // Expected: {'P': 13600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010101; B = 8'b10100000; | Outputs: P=%b | Expected: P=%d",
                 770,
                 
                 P
                 , 
                 
                 13600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101011; B = 8'b01001000; // Expected: {'P': 12312}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101011; B = 8'b01001000; | Outputs: P=%b | Expected: P=%d",
                 771,
                 
                 P
                 , 
                 
                 12312
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000011; B = 8'b10011110; // Expected: {'P': 10586}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000011; B = 8'b10011110; | Outputs: P=%b | Expected: P=%d",
                 772,
                 
                 P
                 , 
                 
                 10586
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001000; B = 8'b11011110; // Expected: {'P': 15984}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001000; B = 8'b11011110; | Outputs: P=%b | Expected: P=%d",
                 773,
                 
                 P
                 , 
                 
                 15984
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001011; B = 8'b00110001; // Expected: {'P': 6811}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001011; B = 8'b00110001; | Outputs: P=%b | Expected: P=%d",
                 774,
                 
                 P
                 , 
                 
                 6811
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100101; B = 8'b01011100; // Expected: {'P': 21068}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100101; B = 8'b01011100; | Outputs: P=%b | Expected: P=%d",
                 775,
                 
                 P
                 , 
                 
                 21068
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111100; B = 8'b11111010; // Expected: {'P': 47000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111100; B = 8'b11111010; | Outputs: P=%b | Expected: P=%d",
                 776,
                 
                 P
                 , 
                 
                 47000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010101; B = 8'b11110111; // Expected: {'P': 5187}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010101; B = 8'b11110111; | Outputs: P=%b | Expected: P=%d",
                 777,
                 
                 P
                 , 
                 
                 5187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001000; B = 8'b00010000; // Expected: {'P': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001000; B = 8'b00010000; | Outputs: P=%b | Expected: P=%d",
                 778,
                 
                 P
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011111; B = 8'b00011001; // Expected: {'P': 775}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011111; B = 8'b00011001; | Outputs: P=%b | Expected: P=%d",
                 779,
                 
                 P
                 , 
                 
                 775
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101101; B = 8'b11101111; // Expected: {'P': 41347}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101101; B = 8'b11101111; | Outputs: P=%b | Expected: P=%d",
                 780,
                 
                 P
                 , 
                 
                 41347
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001000; B = 8'b11001111; // Expected: {'P': 14904}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001000; B = 8'b11001111; | Outputs: P=%b | Expected: P=%d",
                 781,
                 
                 P
                 , 
                 
                 14904
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011111; B = 8'b01110111; // Expected: {'P': 18921}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011111; B = 8'b01110111; | Outputs: P=%b | Expected: P=%d",
                 782,
                 
                 P
                 , 
                 
                 18921
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110110; B = 8'b00001100; // Expected: {'P': 1416}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110110; B = 8'b00001100; | Outputs: P=%b | Expected: P=%d",
                 783,
                 
                 P
                 , 
                 
                 1416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011110; B = 8'b11100010; // Expected: {'P': 50172}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011110; B = 8'b11100010; | Outputs: P=%b | Expected: P=%d",
                 784,
                 
                 P
                 , 
                 
                 50172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000101; B = 8'b01111011; // Expected: {'P': 8487}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000101; B = 8'b01111011; | Outputs: P=%b | Expected: P=%d",
                 785,
                 
                 P
                 , 
                 
                 8487
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110100; B = 8'b01110100; // Expected: {'P': 6032}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110100; B = 8'b01110100; | Outputs: P=%b | Expected: P=%d",
                 786,
                 
                 P
                 , 
                 
                 6032
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010110; B = 8'b00100110; // Expected: {'P': 3268}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010110; B = 8'b00100110; | Outputs: P=%b | Expected: P=%d",
                 787,
                 
                 P
                 , 
                 
                 3268
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101011; B = 8'b11110110; // Expected: {'P': 42066}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101011; B = 8'b11110110; | Outputs: P=%b | Expected: P=%d",
                 788,
                 
                 P
                 , 
                 
                 42066
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110101; B = 8'b01000100; // Expected: {'P': 16660}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110101; B = 8'b01000100; | Outputs: P=%b | Expected: P=%d",
                 789,
                 
                 P
                 , 
                 
                 16660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011101; B = 8'b11010001; // Expected: {'P': 32813}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011101; B = 8'b11010001; | Outputs: P=%b | Expected: P=%d",
                 790,
                 
                 P
                 , 
                 
                 32813
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000000; B = 8'b01100011; // Expected: {'P': 6336}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000000; B = 8'b01100011; | Outputs: P=%b | Expected: P=%d",
                 791,
                 
                 P
                 , 
                 
                 6336
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101000; B = 8'b00101000; // Expected: {'P': 1600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101000; B = 8'b00101000; | Outputs: P=%b | Expected: P=%d",
                 792,
                 
                 P
                 , 
                 
                 1600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100110; B = 8'b01011011; // Expected: {'P': 15106}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100110; B = 8'b01011011; | Outputs: P=%b | Expected: P=%d",
                 793,
                 
                 P
                 , 
                 
                 15106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010111; B = 8'b10011001; // Expected: {'P': 3519}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010111; B = 8'b10011001; | Outputs: P=%b | Expected: P=%d",
                 794,
                 
                 P
                 , 
                 
                 3519
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000110; B = 8'b00011101; // Expected: {'P': 174}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000110; B = 8'b00011101; | Outputs: P=%b | Expected: P=%d",
                 795,
                 
                 P
                 , 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110101; B = 8'b10111101; // Expected: {'P': 22113}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110101; B = 8'b10111101; | Outputs: P=%b | Expected: P=%d",
                 796,
                 
                 P
                 , 
                 
                 22113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000011; B = 8'b11000111; // Expected: {'P': 13333}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000011; B = 8'b11000111; | Outputs: P=%b | Expected: P=%d",
                 797,
                 
                 P
                 , 
                 
                 13333
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101011; B = 8'b11101100; // Expected: {'P': 55460}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101011; B = 8'b11101100; | Outputs: P=%b | Expected: P=%d",
                 798,
                 
                 P
                 , 
                 
                 55460
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000110; B = 8'b10011100; // Expected: {'P': 20904}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000110; B = 8'b10011100; | Outputs: P=%b | Expected: P=%d",
                 799,
                 
                 P
                 , 
                 
                 20904
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001001; B = 8'b10110100; // Expected: {'P': 24660}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001001; B = 8'b10110100; | Outputs: P=%b | Expected: P=%d",
                 800,
                 
                 P
                 , 
                 
                 24660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101001; B = 8'b10010100; // Expected: {'P': 15540}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101001; B = 8'b10010100; | Outputs: P=%b | Expected: P=%d",
                 801,
                 
                 P
                 , 
                 
                 15540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011011; B = 8'b10111100; // Expected: {'P': 5076}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011011; B = 8'b10111100; | Outputs: P=%b | Expected: P=%d",
                 802,
                 
                 P
                 , 
                 
                 5076
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000110; B = 8'b10000011; // Expected: {'P': 9170}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000110; B = 8'b10000011; | Outputs: P=%b | Expected: P=%d",
                 803,
                 
                 P
                 , 
                 
                 9170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001110; B = 8'b00000101; // Expected: {'P': 390}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001110; B = 8'b00000101; | Outputs: P=%b | Expected: P=%d",
                 804,
                 
                 P
                 , 
                 
                 390
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010011; B = 8'b10001011; // Expected: {'P': 11537}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010011; B = 8'b10001011; | Outputs: P=%b | Expected: P=%d",
                 805,
                 
                 P
                 , 
                 
                 11537
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010110; B = 8'b00010011; // Expected: {'P': 2850}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010110; B = 8'b00010011; | Outputs: P=%b | Expected: P=%d",
                 806,
                 
                 P
                 , 
                 
                 2850
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001101; B = 8'b10111000; // Expected: {'P': 2392}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001101; B = 8'b10111000; | Outputs: P=%b | Expected: P=%d",
                 807,
                 
                 P
                 , 
                 
                 2392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101010; B = 8'b01000111; // Expected: {'P': 12070}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101010; B = 8'b01000111; | Outputs: P=%b | Expected: P=%d",
                 808,
                 
                 P
                 , 
                 
                 12070
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100011; B = 8'b11111111; // Expected: {'P': 25245}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100011; B = 8'b11111111; | Outputs: P=%b | Expected: P=%d",
                 809,
                 
                 P
                 , 
                 
                 25245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101111; B = 8'b11001011; // Expected: {'P': 48517}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101111; B = 8'b11001011; | Outputs: P=%b | Expected: P=%d",
                 810,
                 
                 P
                 , 
                 
                 48517
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100110; B = 8'b11101111; // Expected: {'P': 54970}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100110; B = 8'b11101111; | Outputs: P=%b | Expected: P=%d",
                 811,
                 
                 P
                 , 
                 
                 54970
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010111; B = 8'b00000011; // Expected: {'P': 453}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010111; B = 8'b00000011; | Outputs: P=%b | Expected: P=%d",
                 812,
                 
                 P
                 , 
                 
                 453
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001101; B = 8'b11011101; // Expected: {'P': 2873}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001101; B = 8'b11011101; | Outputs: P=%b | Expected: P=%d",
                 813,
                 
                 P
                 , 
                 
                 2873
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111000; B = 8'b00011011; // Expected: {'P': 3240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111000; B = 8'b00011011; | Outputs: P=%b | Expected: P=%d",
                 814,
                 
                 P
                 , 
                 
                 3240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100111; B = 8'b10000100; // Expected: {'P': 22044}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100111; B = 8'b10000100; | Outputs: P=%b | Expected: P=%d",
                 815,
                 
                 P
                 , 
                 
                 22044
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000001; B = 8'b00101001; // Expected: {'P': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000001; B = 8'b00101001; | Outputs: P=%b | Expected: P=%d",
                 816,
                 
                 P
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011000; B = 8'b10100111; // Expected: {'P': 36072}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011000; B = 8'b10100111; | Outputs: P=%b | Expected: P=%d",
                 817,
                 
                 P
                 , 
                 
                 36072
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000001; B = 8'b00011111; // Expected: {'P': 2015}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000001; B = 8'b00011111; | Outputs: P=%b | Expected: P=%d",
                 818,
                 
                 P
                 , 
                 
                 2015
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100110; B = 8'b10001101; // Expected: {'P': 32430}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100110; B = 8'b10001101; | Outputs: P=%b | Expected: P=%d",
                 819,
                 
                 P
                 , 
                 
                 32430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001011; B = 8'b11000010; // Expected: {'P': 2134}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001011; B = 8'b11000010; | Outputs: P=%b | Expected: P=%d",
                 820,
                 
                 P
                 , 
                 
                 2134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111111; B = 8'b10011110; // Expected: {'P': 9954}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111111; B = 8'b10011110; | Outputs: P=%b | Expected: P=%d",
                 821,
                 
                 P
                 , 
                 
                 9954
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101010; B = 8'b01010000; // Expected: {'P': 3360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101010; B = 8'b01010000; | Outputs: P=%b | Expected: P=%d",
                 822,
                 
                 P
                 , 
                 
                 3360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011000; B = 8'b01011001; // Expected: {'P': 13528}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011000; B = 8'b01011001; | Outputs: P=%b | Expected: P=%d",
                 823,
                 
                 P
                 , 
                 
                 13528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110000; B = 8'b11110010; // Expected: {'P': 42592}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110000; B = 8'b11110010; | Outputs: P=%b | Expected: P=%d",
                 824,
                 
                 P
                 , 
                 
                 42592
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000101; B = 8'b00011101; // Expected: {'P': 145}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000101; B = 8'b00011101; | Outputs: P=%b | Expected: P=%d",
                 825,
                 
                 P
                 , 
                 
                 145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000101; B = 8'b01000011; // Expected: {'P': 13199}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000101; B = 8'b01000011; | Outputs: P=%b | Expected: P=%d",
                 826,
                 
                 P
                 , 
                 
                 13199
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000110; B = 8'b00000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000110; B = 8'b00000000; | Outputs: P=%b | Expected: P=%d",
                 827,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001000; B = 8'b01110100; // Expected: {'P': 928}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001000; B = 8'b01110100; | Outputs: P=%b | Expected: P=%d",
                 828,
                 
                 P
                 , 
                 
                 928
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110010; B = 8'b10001011; // Expected: {'P': 24742}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110010; B = 8'b10001011; | Outputs: P=%b | Expected: P=%d",
                 829,
                 
                 P
                 , 
                 
                 24742
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101001; B = 8'b01101111; // Expected: {'P': 11655}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101001; B = 8'b01101111; | Outputs: P=%b | Expected: P=%d",
                 830,
                 
                 P
                 , 
                 
                 11655
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000100; B = 8'b01000111; // Expected: {'P': 9372}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000100; B = 8'b01000111; | Outputs: P=%b | Expected: P=%d",
                 831,
                 
                 P
                 , 
                 
                 9372
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010100; B = 8'b10001001; // Expected: {'P': 29044}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010100; B = 8'b10001001; | Outputs: P=%b | Expected: P=%d",
                 832,
                 
                 P
                 , 
                 
                 29044
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001001; B = 8'b11110010; // Expected: {'P': 2178}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001001; B = 8'b11110010; | Outputs: P=%b | Expected: P=%d",
                 833,
                 
                 P
                 , 
                 
                 2178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101100; B = 8'b10111011; // Expected: {'P': 20196}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101100; B = 8'b10111011; | Outputs: P=%b | Expected: P=%d",
                 834,
                 
                 P
                 , 
                 
                 20196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000000; B = 8'b00011011; // Expected: {'P': 5184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000000; B = 8'b00011011; | Outputs: P=%b | Expected: P=%d",
                 835,
                 
                 P
                 , 
                 
                 5184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100100; B = 8'b11110100; // Expected: {'P': 40016}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100100; B = 8'b11110100; | Outputs: P=%b | Expected: P=%d",
                 836,
                 
                 P
                 , 
                 
                 40016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001010; B = 8'b01000001; // Expected: {'P': 650}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001010; B = 8'b01000001; | Outputs: P=%b | Expected: P=%d",
                 837,
                 
                 P
                 , 
                 
                 650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011001; B = 8'b10110101; // Expected: {'P': 27693}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011001; B = 8'b10110101; | Outputs: P=%b | Expected: P=%d",
                 838,
                 
                 P
                 , 
                 
                 27693
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010011; B = 8'b00010101; // Expected: {'P': 3087}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010011; B = 8'b00010101; | Outputs: P=%b | Expected: P=%d",
                 839,
                 
                 P
                 , 
                 
                 3087
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011110; B = 8'b11011100; // Expected: {'P': 20680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011110; B = 8'b11011100; | Outputs: P=%b | Expected: P=%d",
                 840,
                 
                 P
                 , 
                 
                 20680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001110; B = 8'b00110101; // Expected: {'P': 10918}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001110; B = 8'b00110101; | Outputs: P=%b | Expected: P=%d",
                 841,
                 
                 P
                 , 
                 
                 10918
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001001; B = 8'b01111011; // Expected: {'P': 16851}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001001; B = 8'b01111011; | Outputs: P=%b | Expected: P=%d",
                 842,
                 
                 P
                 , 
                 
                 16851
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001011; B = 8'b00101100; // Expected: {'P': 6116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001011; B = 8'b00101100; | Outputs: P=%b | Expected: P=%d",
                 843,
                 
                 P
                 , 
                 
                 6116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110111; B = 8'b01101110; // Expected: {'P': 13090}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110111; B = 8'b01101110; | Outputs: P=%b | Expected: P=%d",
                 844,
                 
                 P
                 , 
                 
                 13090
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110101; B = 8'b10100011; // Expected: {'P': 29503}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110101; B = 8'b10100011; | Outputs: P=%b | Expected: P=%d",
                 845,
                 
                 P
                 , 
                 
                 29503
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111110; B = 8'b11101001; // Expected: {'P': 59182}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111110; B = 8'b11101001; | Outputs: P=%b | Expected: P=%d",
                 846,
                 
                 P
                 , 
                 
                 59182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011010; B = 8'b00010101; // Expected: {'P': 546}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011010; B = 8'b00010101; | Outputs: P=%b | Expected: P=%d",
                 847,
                 
                 P
                 , 
                 
                 546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010001; B = 8'b10001010; // Expected: {'P': 28842}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010001; B = 8'b10001010; | Outputs: P=%b | Expected: P=%d",
                 848,
                 
                 P
                 , 
                 
                 28842
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101111; B = 8'b00001011; // Expected: {'P': 517}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101111; B = 8'b00001011; | Outputs: P=%b | Expected: P=%d",
                 849,
                 
                 P
                 , 
                 
                 517
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101000; B = 8'b01011111; // Expected: {'P': 15960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101000; B = 8'b01011111; | Outputs: P=%b | Expected: P=%d",
                 850,
                 
                 P
                 , 
                 
                 15960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101010; B = 8'b01100000; // Expected: {'P': 10176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101010; B = 8'b01100000; | Outputs: P=%b | Expected: P=%d",
                 851,
                 
                 P
                 , 
                 
                 10176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001010; B = 8'b01011001; // Expected: {'P': 890}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001010; B = 8'b01011001; | Outputs: P=%b | Expected: P=%d",
                 852,
                 
                 P
                 , 
                 
                 890
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010110; B = 8'b01001010; // Expected: {'P': 15836}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010110; B = 8'b01001010; | Outputs: P=%b | Expected: P=%d",
                 853,
                 
                 P
                 , 
                 
                 15836
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101100; B = 8'b00011101; // Expected: {'P': 6844}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101100; B = 8'b00011101; | Outputs: P=%b | Expected: P=%d",
                 854,
                 
                 P
                 , 
                 
                 6844
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101100; B = 8'b01010010; // Expected: {'P': 14104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101100; B = 8'b01010010; | Outputs: P=%b | Expected: P=%d",
                 855,
                 
                 P
                 , 
                 
                 14104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001000; B = 8'b01010000; // Expected: {'P': 10880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001000; B = 8'b01010000; | Outputs: P=%b | Expected: P=%d",
                 856,
                 
                 P
                 , 
                 
                 10880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010100; B = 8'b00110110; // Expected: {'P': 11448}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010100; B = 8'b00110110; | Outputs: P=%b | Expected: P=%d",
                 857,
                 
                 P
                 , 
                 
                 11448
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100111; B = 8'b01110110; // Expected: {'P': 12154}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100111; B = 8'b01110110; | Outputs: P=%b | Expected: P=%d",
                 858,
                 
                 P
                 , 
                 
                 12154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010111; B = 8'b00001110; // Expected: {'P': 322}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010111; B = 8'b00001110; | Outputs: P=%b | Expected: P=%d",
                 859,
                 
                 P
                 , 
                 
                 322
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010010; B = 8'b11110101; // Expected: {'P': 51450}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010010; B = 8'b11110101; | Outputs: P=%b | Expected: P=%d",
                 860,
                 
                 P
                 , 
                 
                 51450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110000; B = 8'b10011000; // Expected: {'P': 7296}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110000; B = 8'b10011000; | Outputs: P=%b | Expected: P=%d",
                 861,
                 
                 P
                 , 
                 
                 7296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101111; B = 8'b01011100; // Expected: {'P': 21988}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101111; B = 8'b01011100; | Outputs: P=%b | Expected: P=%d",
                 862,
                 
                 P
                 , 
                 
                 21988
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000100; B = 8'b00011111; // Expected: {'P': 4092}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000100; B = 8'b00011111; | Outputs: P=%b | Expected: P=%d",
                 863,
                 
                 P
                 , 
                 
                 4092
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110110; B = 8'b10110011; // Expected: {'P': 32578}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110110; B = 8'b10110011; | Outputs: P=%b | Expected: P=%d",
                 864,
                 
                 P
                 , 
                 
                 32578
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000101; B = 8'b11011011; // Expected: {'P': 43143}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000101; B = 8'b11011011; | Outputs: P=%b | Expected: P=%d",
                 865,
                 
                 P
                 , 
                 
                 43143
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011100; B = 8'b01111010; // Expected: {'P': 11224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011100; B = 8'b01111010; | Outputs: P=%b | Expected: P=%d",
                 866,
                 
                 P
                 , 
                 
                 11224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011110; B = 8'b10000110; // Expected: {'P': 21172}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011110; B = 8'b10000110; | Outputs: P=%b | Expected: P=%d",
                 867,
                 
                 P
                 , 
                 
                 21172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010111; B = 8'b00001010; // Expected: {'P': 2150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010111; B = 8'b00001010; | Outputs: P=%b | Expected: P=%d",
                 868,
                 
                 P
                 , 
                 
                 2150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000001; B = 8'b01001011; // Expected: {'P': 9675}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000001; B = 8'b01001011; | Outputs: P=%b | Expected: P=%d",
                 869,
                 
                 P
                 , 
                 
                 9675
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101000; B = 8'b11101000; // Expected: {'P': 9280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101000; B = 8'b11101000; | Outputs: P=%b | Expected: P=%d",
                 870,
                 
                 P
                 , 
                 
                 9280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001010; B = 8'b01111001; // Expected: {'P': 1210}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001010; B = 8'b01111001; | Outputs: P=%b | Expected: P=%d",
                 871,
                 
                 P
                 , 
                 
                 1210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001010; B = 8'b10110101; // Expected: {'P': 1810}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001010; B = 8'b10110101; | Outputs: P=%b | Expected: P=%d",
                 872,
                 
                 P
                 , 
                 
                 1810
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010010; B = 8'b01101100; // Expected: {'P': 22680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010010; B = 8'b01101100; | Outputs: P=%b | Expected: P=%d",
                 873,
                 
                 P
                 , 
                 
                 22680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110111; B = 8'b10010010; // Expected: {'P': 26718}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110111; B = 8'b10010010; | Outputs: P=%b | Expected: P=%d",
                 874,
                 
                 P
                 , 
                 
                 26718
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110100; B = 8'b10110100; // Expected: {'P': 20880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110100; B = 8'b10110100; | Outputs: P=%b | Expected: P=%d",
                 875,
                 
                 P
                 , 
                 
                 20880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111000; B = 8'b11100010; // Expected: {'P': 27120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111000; B = 8'b11100010; | Outputs: P=%b | Expected: P=%d",
                 876,
                 
                 P
                 , 
                 
                 27120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111010; B = 8'b11101111; // Expected: {'P': 44454}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111010; B = 8'b11101111; | Outputs: P=%b | Expected: P=%d",
                 877,
                 
                 P
                 , 
                 
                 44454
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111111; B = 8'b01011100; // Expected: {'P': 5796}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111111; B = 8'b01011100; | Outputs: P=%b | Expected: P=%d",
                 878,
                 
                 P
                 , 
                 
                 5796
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000101; B = 8'b00100100; // Expected: {'P': 7092}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000101; B = 8'b00100100; | Outputs: P=%b | Expected: P=%d",
                 879,
                 
                 P
                 , 
                 
                 7092
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011000; B = 8'b11001100; // Expected: {'P': 17952}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011000; B = 8'b11001100; | Outputs: P=%b | Expected: P=%d",
                 880,
                 
                 P
                 , 
                 
                 17952
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101010; B = 8'b00000110; // Expected: {'P': 1404}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101010; B = 8'b00000110; | Outputs: P=%b | Expected: P=%d",
                 881,
                 
                 P
                 , 
                 
                 1404
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001011; B = 8'b11001101; // Expected: {'P': 15375}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001011; B = 8'b11001101; | Outputs: P=%b | Expected: P=%d",
                 882,
                 
                 P
                 , 
                 
                 15375
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111100; B = 8'b10011101; // Expected: {'P': 39564}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111100; B = 8'b10011101; | Outputs: P=%b | Expected: P=%d",
                 883,
                 
                 P
                 , 
                 
                 39564
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110011; B = 8'b01100001; // Expected: {'P': 4947}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110011; B = 8'b01100001; | Outputs: P=%b | Expected: P=%d",
                 884,
                 
                 P
                 , 
                 
                 4947
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000011; B = 8'b10111111; // Expected: {'P': 573}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000011; B = 8'b10111111; | Outputs: P=%b | Expected: P=%d",
                 885,
                 
                 P
                 , 
                 
                 573
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100101; B = 8'b11111010; // Expected: {'P': 57250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100101; B = 8'b11111010; | Outputs: P=%b | Expected: P=%d",
                 886,
                 
                 P
                 , 
                 
                 57250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000011; B = 8'b11010110; // Expected: {'P': 28034}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000011; B = 8'b11010110; | Outputs: P=%b | Expected: P=%d",
                 887,
                 
                 P
                 , 
                 
                 28034
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110111; B = 8'b10000000; // Expected: {'P': 23424}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110111; B = 8'b10000000; | Outputs: P=%b | Expected: P=%d",
                 888,
                 
                 P
                 , 
                 
                 23424
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010110; B = 8'b10111001; // Expected: {'P': 4070}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010110; B = 8'b10111001; | Outputs: P=%b | Expected: P=%d",
                 889,
                 
                 P
                 , 
                 
                 4070
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100110; B = 8'b11011111; // Expected: {'P': 51290}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100110; B = 8'b11011111; | Outputs: P=%b | Expected: P=%d",
                 890,
                 
                 P
                 , 
                 
                 51290
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101000; B = 8'b00010001; // Expected: {'P': 680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101000; B = 8'b00010001; | Outputs: P=%b | Expected: P=%d",
                 891,
                 
                 P
                 , 
                 
                 680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110111; B = 8'b10010100; // Expected: {'P': 36556}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110111; B = 8'b10010100; | Outputs: P=%b | Expected: P=%d",
                 892,
                 
                 P
                 , 
                 
                 36556
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101110; B = 8'b01111101; // Expected: {'P': 13750}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101110; B = 8'b01111101; | Outputs: P=%b | Expected: P=%d",
                 893,
                 
                 P
                 , 
                 
                 13750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100011; B = 8'b00001111; // Expected: {'P': 3405}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100011; B = 8'b00001111; | Outputs: P=%b | Expected: P=%d",
                 894,
                 
                 P
                 , 
                 
                 3405
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101100; B = 8'b00100000; // Expected: {'P': 5504}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101100; B = 8'b00100000; | Outputs: P=%b | Expected: P=%d",
                 895,
                 
                 P
                 , 
                 
                 5504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001001; B = 8'b00000001; // Expected: {'P': 73}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001001; B = 8'b00000001; | Outputs: P=%b | Expected: P=%d",
                 896,
                 
                 P
                 , 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010110; B = 8'b00001100; // Expected: {'P': 1800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010110; B = 8'b00001100; | Outputs: P=%b | Expected: P=%d",
                 897,
                 
                 P
                 , 
                 
                 1800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000101; B = 8'b11101001; // Expected: {'P': 30989}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000101; B = 8'b11101001; | Outputs: P=%b | Expected: P=%d",
                 898,
                 
                 P
                 , 
                 
                 30989
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000111; B = 8'b10011110; // Expected: {'P': 21330}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000111; B = 8'b10011110; | Outputs: P=%b | Expected: P=%d",
                 899,
                 
                 P
                 , 
                 
                 21330
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001011; B = 8'b00001100; // Expected: {'P': 900}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001011; B = 8'b00001100; | Outputs: P=%b | Expected: P=%d",
                 900,
                 
                 P
                 , 
                 
                 900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001000; B = 8'b10111001; // Expected: {'P': 37000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001000; B = 8'b10111001; | Outputs: P=%b | Expected: P=%d",
                 901,
                 
                 P
                 , 
                 
                 37000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100110; B = 8'b11111011; // Expected: {'P': 25602}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100110; B = 8'b11111011; | Outputs: P=%b | Expected: P=%d",
                 902,
                 
                 P
                 , 
                 
                 25602
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010011; B = 8'b00000111; // Expected: {'P': 1477}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010011; B = 8'b00000111; | Outputs: P=%b | Expected: P=%d",
                 903,
                 
                 P
                 , 
                 
                 1477
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101011; B = 8'b00000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101011; B = 8'b00000000; | Outputs: P=%b | Expected: P=%d",
                 904,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101110; B = 8'b11011010; // Expected: {'P': 51884}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101110; B = 8'b11011010; | Outputs: P=%b | Expected: P=%d",
                 905,
                 
                 P
                 , 
                 
                 51884
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011100; B = 8'b01100000; // Expected: {'P': 14976}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011100; B = 8'b01100000; | Outputs: P=%b | Expected: P=%d",
                 906,
                 
                 P
                 , 
                 
                 14976
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100111; B = 8'b10101001; // Expected: {'P': 39039}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100111; B = 8'b10101001; | Outputs: P=%b | Expected: P=%d",
                 907,
                 
                 P
                 , 
                 
                 39039
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101101; B = 8'b00000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101101; B = 8'b00000000; | Outputs: P=%b | Expected: P=%d",
                 908,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010001; B = 8'b11010001; // Expected: {'P': 30305}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010001; B = 8'b11010001; | Outputs: P=%b | Expected: P=%d",
                 909,
                 
                 P
                 , 
                 
                 30305
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001100; B = 8'b10101010; // Expected: {'P': 23800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001100; B = 8'b10101010; | Outputs: P=%b | Expected: P=%d",
                 910,
                 
                 P
                 , 
                 
                 23800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011001; B = 8'b10000001; // Expected: {'P': 3225}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011001; B = 8'b10000001; | Outputs: P=%b | Expected: P=%d",
                 911,
                 
                 P
                 , 
                 
                 3225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110110; B = 8'b10111110; // Expected: {'P': 22420}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110110; B = 8'b10111110; | Outputs: P=%b | Expected: P=%d",
                 912,
                 
                 P
                 , 
                 
                 22420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011101; B = 8'b00110010; // Expected: {'P': 7850}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011101; B = 8'b00110010; | Outputs: P=%b | Expected: P=%d",
                 913,
                 
                 P
                 , 
                 
                 7850
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010000; B = 8'b01001110; // Expected: {'P': 6240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010000; B = 8'b01001110; | Outputs: P=%b | Expected: P=%d",
                 914,
                 
                 P
                 , 
                 
                 6240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011000; B = 8'b10111111; // Expected: {'P': 29032}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011000; B = 8'b10111111; | Outputs: P=%b | Expected: P=%d",
                 915,
                 
                 P
                 , 
                 
                 29032
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101110; B = 8'b01001111; // Expected: {'P': 3634}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101110; B = 8'b01001111; | Outputs: P=%b | Expected: P=%d",
                 916,
                 
                 P
                 , 
                 
                 3634
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010100; B = 8'b11101000; // Expected: {'P': 34336}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010100; B = 8'b11101000; | Outputs: P=%b | Expected: P=%d",
                 917,
                 
                 P
                 , 
                 
                 34336
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111000; B = 8'b11010110; // Expected: {'P': 39376}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111000; B = 8'b11010110; | Outputs: P=%b | Expected: P=%d",
                 918,
                 
                 P
                 , 
                 
                 39376
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000011; B = 8'b10011000; // Expected: {'P': 456}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000011; B = 8'b10011000; | Outputs: P=%b | Expected: P=%d",
                 919,
                 
                 P
                 , 
                 
                 456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100010; B = 8'b11001001; // Expected: {'P': 45426}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100010; B = 8'b11001001; | Outputs: P=%b | Expected: P=%d",
                 920,
                 
                 P
                 , 
                 
                 45426
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001101; B = 8'b10001100; // Expected: {'P': 1820}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001101; B = 8'b10001100; | Outputs: P=%b | Expected: P=%d",
                 921,
                 
                 P
                 , 
                 
                 1820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101100; B = 8'b01101010; // Expected: {'P': 4664}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101100; B = 8'b01101010; | Outputs: P=%b | Expected: P=%d",
                 922,
                 
                 P
                 , 
                 
                 4664
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111110; B = 8'b11101101; // Expected: {'P': 60198}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111110; B = 8'b11101101; | Outputs: P=%b | Expected: P=%d",
                 923,
                 
                 P
                 , 
                 
                 60198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101001; B = 8'b11110000; // Expected: {'P': 55920}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101001; B = 8'b11110000; | Outputs: P=%b | Expected: P=%d",
                 924,
                 
                 P
                 , 
                 
                 55920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010000; B = 8'b00100101; // Expected: {'P': 7696}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010000; B = 8'b00100101; | Outputs: P=%b | Expected: P=%d",
                 925,
                 
                 P
                 , 
                 
                 7696
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010001; B = 8'b00110110; // Expected: {'P': 918}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010001; B = 8'b00110110; | Outputs: P=%b | Expected: P=%d",
                 926,
                 
                 P
                 , 
                 
                 918
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011001; B = 8'b11100111; // Expected: {'P': 20559}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011001; B = 8'b11100111; | Outputs: P=%b | Expected: P=%d",
                 927,
                 
                 P
                 , 
                 
                 20559
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001100; B = 8'b10110110; // Expected: {'P': 2184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001100; B = 8'b10110110; | Outputs: P=%b | Expected: P=%d",
                 928,
                 
                 P
                 , 
                 
                 2184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101000; B = 8'b11011000; // Expected: {'P': 36288}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101000; B = 8'b11011000; | Outputs: P=%b | Expected: P=%d",
                 929,
                 
                 P
                 , 
                 
                 36288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110111; B = 8'b10011111; // Expected: {'P': 18921}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110111; B = 8'b10011111; | Outputs: P=%b | Expected: P=%d",
                 930,
                 
                 P
                 , 
                 
                 18921
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110101; B = 8'b01111100; // Expected: {'P': 6572}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110101; B = 8'b01111100; | Outputs: P=%b | Expected: P=%d",
                 931,
                 
                 P
                 , 
                 
                 6572
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101000; B = 8'b00011111; // Expected: {'P': 5208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101000; B = 8'b00011111; | Outputs: P=%b | Expected: P=%d",
                 932,
                 
                 P
                 , 
                 
                 5208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111011; B = 8'b00010100; // Expected: {'P': 2460}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111011; B = 8'b00010100; | Outputs: P=%b | Expected: P=%d",
                 933,
                 
                 P
                 , 
                 
                 2460
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000011; B = 8'b01110110; // Expected: {'P': 23010}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000011; B = 8'b01110110; | Outputs: P=%b | Expected: P=%d",
                 934,
                 
                 P
                 , 
                 
                 23010
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010010; B = 8'b00101100; // Expected: {'P': 792}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010010; B = 8'b00101100; | Outputs: P=%b | Expected: P=%d",
                 935,
                 
                 P
                 , 
                 
                 792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100000; B = 8'b01011001; // Expected: {'P': 8544}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100000; B = 8'b01011001; | Outputs: P=%b | Expected: P=%d",
                 936,
                 
                 P
                 , 
                 
                 8544
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001011; B = 8'b11001001; // Expected: {'P': 27939}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001011; B = 8'b11001001; | Outputs: P=%b | Expected: P=%d",
                 937,
                 
                 P
                 , 
                 
                 27939
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100001; B = 8'b11110010; // Expected: {'P': 23474}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100001; B = 8'b11110010; | Outputs: P=%b | Expected: P=%d",
                 938,
                 
                 P
                 , 
                 
                 23474
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001011; B = 8'b00110111; // Expected: {'P': 11165}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001011; B = 8'b00110111; | Outputs: P=%b | Expected: P=%d",
                 939,
                 
                 P
                 , 
                 
                 11165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111100; B = 8'b01101010; // Expected: {'P': 13144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111100; B = 8'b01101010; | Outputs: P=%b | Expected: P=%d",
                 940,
                 
                 P
                 , 
                 
                 13144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110011; B = 8'b10000110; // Expected: {'P': 32562}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110011; B = 8'b10000110; | Outputs: P=%b | Expected: P=%d",
                 941,
                 
                 P
                 , 
                 
                 32562
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111011; B = 8'b01000000; // Expected: {'P': 16064}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111011; B = 8'b01000000; | Outputs: P=%b | Expected: P=%d",
                 942,
                 
                 P
                 , 
                 
                 16064
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101110; B = 8'b11100101; // Expected: {'P': 39846}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101110; B = 8'b11100101; | Outputs: P=%b | Expected: P=%d",
                 943,
                 
                 P
                 , 
                 
                 39846
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101010; B = 8'b01011111; // Expected: {'P': 3990}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101010; B = 8'b01011111; | Outputs: P=%b | Expected: P=%d",
                 944,
                 
                 P
                 , 
                 
                 3990
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000000; B = 8'b01011100; // Expected: {'P': 11776}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000000; B = 8'b01011100; | Outputs: P=%b | Expected: P=%d",
                 945,
                 
                 P
                 , 
                 
                 11776
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000001; B = 8'b00100111; // Expected: {'P': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000001; B = 8'b00100111; | Outputs: P=%b | Expected: P=%d",
                 946,
                 
                 P
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011110; B = 8'b00110110; // Expected: {'P': 5076}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011110; B = 8'b00110110; | Outputs: P=%b | Expected: P=%d",
                 947,
                 
                 P
                 , 
                 
                 5076
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101001; B = 8'b00001100; // Expected: {'P': 492}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101001; B = 8'b00001100; | Outputs: P=%b | Expected: P=%d",
                 948,
                 
                 P
                 , 
                 
                 492
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101011; B = 8'b11011011; // Expected: {'P': 9417}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101011; B = 8'b11011011; | Outputs: P=%b | Expected: P=%d",
                 949,
                 
                 P
                 , 
                 
                 9417
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110011; B = 8'b01000010; // Expected: {'P': 11814}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110011; B = 8'b01000010; | Outputs: P=%b | Expected: P=%d",
                 950,
                 
                 P
                 , 
                 
                 11814
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011101; B = 8'b00110101; // Expected: {'P': 1537}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011101; B = 8'b00110101; | Outputs: P=%b | Expected: P=%d",
                 951,
                 
                 P
                 , 
                 
                 1537
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011010; B = 8'b01011000; // Expected: {'P': 19184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011010; B = 8'b01011000; | Outputs: P=%b | Expected: P=%d",
                 952,
                 
                 P
                 , 
                 
                 19184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100011; B = 8'b10000011; // Expected: {'P': 4585}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100011; B = 8'b10000011; | Outputs: P=%b | Expected: P=%d",
                 953,
                 
                 P
                 , 
                 
                 4585
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001100; B = 8'b01000000; // Expected: {'P': 8960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001100; B = 8'b01000000; | Outputs: P=%b | Expected: P=%d",
                 954,
                 
                 P
                 , 
                 
                 8960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010001; B = 8'b10110110; // Expected: {'P': 14742}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010001; B = 8'b10110110; | Outputs: P=%b | Expected: P=%d",
                 955,
                 
                 P
                 , 
                 
                 14742
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111000; B = 8'b10101110; // Expected: {'P': 32016}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111000; B = 8'b10101110; | Outputs: P=%b | Expected: P=%d",
                 956,
                 
                 P
                 , 
                 
                 32016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101001; B = 8'b10100000; // Expected: {'P': 27040}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101001; B = 8'b10100000; | Outputs: P=%b | Expected: P=%d",
                 957,
                 
                 P
                 , 
                 
                 27040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100100; B = 8'b10010100; // Expected: {'P': 5328}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100100; B = 8'b10010100; | Outputs: P=%b | Expected: P=%d",
                 958,
                 
                 P
                 , 
                 
                 5328
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000101; B = 8'b01010110; // Expected: {'P': 430}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000101; B = 8'b01010110; | Outputs: P=%b | Expected: P=%d",
                 959,
                 
                 P
                 , 
                 
                 430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001100; B = 8'b10001101; // Expected: {'P': 1692}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001100; B = 8'b10001101; | Outputs: P=%b | Expected: P=%d",
                 960,
                 
                 P
                 , 
                 
                 1692
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110011; B = 8'b00011001; // Expected: {'P': 2875}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110011; B = 8'b00011001; | Outputs: P=%b | Expected: P=%d",
                 961,
                 
                 P
                 , 
                 
                 2875
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001101; B = 8'b10100010; // Expected: {'P': 33210}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001101; B = 8'b10100010; | Outputs: P=%b | Expected: P=%d",
                 962,
                 
                 P
                 , 
                 
                 33210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100101; B = 8'b11001000; // Expected: {'P': 7400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100101; B = 8'b11001000; | Outputs: P=%b | Expected: P=%d",
                 963,
                 
                 P
                 , 
                 
                 7400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001110; B = 8'b01011001; // Expected: {'P': 1246}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001110; B = 8'b01011001; | Outputs: P=%b | Expected: P=%d",
                 964,
                 
                 P
                 , 
                 
                 1246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100111; B = 8'b01000000; // Expected: {'P': 2496}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100111; B = 8'b01000000; | Outputs: P=%b | Expected: P=%d",
                 965,
                 
                 P
                 , 
                 
                 2496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100100; B = 8'b00010011; // Expected: {'P': 1900}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100100; B = 8'b00010011; | Outputs: P=%b | Expected: P=%d",
                 966,
                 
                 P
                 , 
                 
                 1900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110010; B = 8'b10000001; // Expected: {'P': 22962}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110010; B = 8'b10000001; | Outputs: P=%b | Expected: P=%d",
                 967,
                 
                 P
                 , 
                 
                 22962
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011011; B = 8'b10110011; // Expected: {'P': 4833}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011011; B = 8'b10110011; | Outputs: P=%b | Expected: P=%d",
                 968,
                 
                 P
                 , 
                 
                 4833
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110101; B = 8'b01011000; // Expected: {'P': 21560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110101; B = 8'b01011000; | Outputs: P=%b | Expected: P=%d",
                 969,
                 
                 P
                 , 
                 
                 21560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011011; B = 8'b00000001; // Expected: {'P': 91}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011011; B = 8'b00000001; | Outputs: P=%b | Expected: P=%d",
                 970,
                 
                 P
                 , 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100111; B = 8'b11000011; // Expected: {'P': 45045}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100111; B = 8'b11000011; | Outputs: P=%b | Expected: P=%d",
                 971,
                 
                 P
                 , 
                 
                 45045
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001111; B = 8'b00001011; // Expected: {'P': 1573}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001111; B = 8'b00001011; | Outputs: P=%b | Expected: P=%d",
                 972,
                 
                 P
                 , 
                 
                 1573
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100110; B = 8'b10010001; // Expected: {'P': 33350}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100110; B = 8'b10010001; | Outputs: P=%b | Expected: P=%d",
                 973,
                 
                 P
                 , 
                 
                 33350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010110; B = 8'b11111110; // Expected: {'P': 38100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010110; B = 8'b11111110; | Outputs: P=%b | Expected: P=%d",
                 974,
                 
                 P
                 , 
                 
                 38100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101111; B = 8'b10010001; // Expected: {'P': 34655}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101111; B = 8'b10010001; | Outputs: P=%b | Expected: P=%d",
                 975,
                 
                 P
                 , 
                 
                 34655
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011000; B = 8'b10011110; // Expected: {'P': 3792}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011000; B = 8'b10011110; | Outputs: P=%b | Expected: P=%d",
                 976,
                 
                 P
                 , 
                 
                 3792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110000; B = 8'b10011111; // Expected: {'P': 17808}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110000; B = 8'b10011111; | Outputs: P=%b | Expected: P=%d",
                 977,
                 
                 P
                 , 
                 
                 17808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110011; B = 8'b10001110; // Expected: {'P': 34506}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110011; B = 8'b10001110; | Outputs: P=%b | Expected: P=%d",
                 978,
                 
                 P
                 , 
                 
                 34506
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000000; B = 8'b11111101; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000000; B = 8'b11111101; | Outputs: P=%b | Expected: P=%d",
                 979,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011010; B = 8'b01010101; // Expected: {'P': 2210}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011010; B = 8'b01010101; | Outputs: P=%b | Expected: P=%d",
                 980,
                 
                 P
                 , 
                 
                 2210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111001; B = 8'b10001000; // Expected: {'P': 33864}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111001; B = 8'b10001000; | Outputs: P=%b | Expected: P=%d",
                 981,
                 
                 P
                 , 
                 
                 33864
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110011; B = 8'b10011100; // Expected: {'P': 17940}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110011; B = 8'b10011100; | Outputs: P=%b | Expected: P=%d",
                 982,
                 
                 P
                 , 
                 
                 17940
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101111; B = 8'b11011001; // Expected: {'P': 24087}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101111; B = 8'b11011001; | Outputs: P=%b | Expected: P=%d",
                 983,
                 
                 P
                 , 
                 
                 24087
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101100; B = 8'b01000100; // Expected: {'P': 11696}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101100; B = 8'b01000100; | Outputs: P=%b | Expected: P=%d",
                 984,
                 
                 P
                 , 
                 
                 11696
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010101; B = 8'b00101110; // Expected: {'P': 9798}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010101; B = 8'b00101110; | Outputs: P=%b | Expected: P=%d",
                 985,
                 
                 P
                 , 
                 
                 9798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110011; B = 8'b01000101; // Expected: {'P': 7935}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110011; B = 8'b01000101; | Outputs: P=%b | Expected: P=%d",
                 986,
                 
                 P
                 , 
                 
                 7935
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101001; B = 8'b10100000; // Expected: {'P': 16800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101001; B = 8'b10100000; | Outputs: P=%b | Expected: P=%d",
                 987,
                 
                 P
                 , 
                 
                 16800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001101; B = 8'b00110000; // Expected: {'P': 9840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001101; B = 8'b00110000; | Outputs: P=%b | Expected: P=%d",
                 988,
                 
                 P
                 , 
                 
                 9840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101011; B = 8'b11001110; // Expected: {'P': 8858}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101011; B = 8'b11001110; | Outputs: P=%b | Expected: P=%d",
                 989,
                 
                 P
                 , 
                 
                 8858
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110100; B = 8'b00010100; // Expected: {'P': 2320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110100; B = 8'b00010100; | Outputs: P=%b | Expected: P=%d",
                 990,
                 
                 P
                 , 
                 
                 2320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010000; B = 8'b01001010; // Expected: {'P': 15392}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010000; B = 8'b01001010; | Outputs: P=%b | Expected: P=%d",
                 991,
                 
                 P
                 , 
                 
                 15392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011111; B = 8'b01001110; // Expected: {'P': 2418}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011111; B = 8'b01001110; | Outputs: P=%b | Expected: P=%d",
                 992,
                 
                 P
                 , 
                 
                 2418
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101101; B = 8'b01100011; // Expected: {'P': 4455}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101101; B = 8'b01100011; | Outputs: P=%b | Expected: P=%d",
                 993,
                 
                 P
                 , 
                 
                 4455
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000011; B = 8'b00100011; // Expected: {'P': 4585}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000011; B = 8'b00100011; | Outputs: P=%b | Expected: P=%d",
                 994,
                 
                 P
                 , 
                 
                 4585
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000001; B = 8'b01010010; // Expected: {'P': 82}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000001; B = 8'b01010010; | Outputs: P=%b | Expected: P=%d",
                 995,
                 
                 P
                 , 
                 
                 82
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101100; B = 8'b11010000; // Expected: {'P': 22464}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101100; B = 8'b11010000; | Outputs: P=%b | Expected: P=%d",
                 996,
                 
                 P
                 , 
                 
                 22464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000101; B = 8'b10100100; // Expected: {'P': 820}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000101; B = 8'b10100100; | Outputs: P=%b | Expected: P=%d",
                 997,
                 
                 P
                 , 
                 
                 820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110001; B = 8'b11111001; // Expected: {'P': 44073}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110001; B = 8'b11111001; | Outputs: P=%b | Expected: P=%d",
                 998,
                 
                 P
                 , 
                 
                 44073
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111101; B = 8'b01110011; // Expected: {'P': 21735}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111101; B = 8'b01110011; | Outputs: P=%b | Expected: P=%d",
                 999,
                 
                 P
                 , 
                 
                 21735
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110001; B = 8'b00100100; // Expected: {'P': 4068}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110001; B = 8'b00100100; | Outputs: P=%b | Expected: P=%d",
                 1000,
                 
                 P
                 , 
                 
                 4068
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111110; B = 8'b11101011; // Expected: {'P': 14570}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111110; B = 8'b11101011; | Outputs: P=%b | Expected: P=%d",
                 1001,
                 
                 P
                 , 
                 
                 14570
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000111; B = 8'b10101110; // Expected: {'P': 23490}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000111; B = 8'b10101110; | Outputs: P=%b | Expected: P=%d",
                 1002,
                 
                 P
                 , 
                 
                 23490
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001111; B = 8'b11110000; // Expected: {'P': 3600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001111; B = 8'b11110000; | Outputs: P=%b | Expected: P=%d",
                 1003,
                 
                 P
                 , 
                 
                 3600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101111; B = 8'b10101100; // Expected: {'P': 30100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101111; B = 8'b10101100; | Outputs: P=%b | Expected: P=%d",
                 1004,
                 
                 P
                 , 
                 
                 30100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101010; B = 8'b10101011; // Expected: {'P': 40014}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101010; B = 8'b10101011; | Outputs: P=%b | Expected: P=%d",
                 1005,
                 
                 P
                 , 
                 
                 40014
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110111; B = 8'b01011110; // Expected: {'P': 11186}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110111; B = 8'b01011110; | Outputs: P=%b | Expected: P=%d",
                 1006,
                 
                 P
                 , 
                 
                 11186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001011; B = 8'b11101111; // Expected: {'P': 33221}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001011; B = 8'b11101111; | Outputs: P=%b | Expected: P=%d",
                 1007,
                 
                 P
                 , 
                 
                 33221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010111; B = 8'b00111000; // Expected: {'P': 8456}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010111; B = 8'b00111000; | Outputs: P=%b | Expected: P=%d",
                 1008,
                 
                 P
                 , 
                 
                 8456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101101; B = 8'b01110011; // Expected: {'P': 5175}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101101; B = 8'b01110011; | Outputs: P=%b | Expected: P=%d",
                 1009,
                 
                 P
                 , 
                 
                 5175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101111; B = 8'b10011101; // Expected: {'P': 7379}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101111; B = 8'b10011101; | Outputs: P=%b | Expected: P=%d",
                 1010,
                 
                 P
                 , 
                 
                 7379
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101001; B = 8'b01100011; // Expected: {'P': 16731}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101001; B = 8'b01100011; | Outputs: P=%b | Expected: P=%d",
                 1011,
                 
                 P
                 , 
                 
                 16731
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111110; B = 8'b10110111; // Expected: {'P': 11346}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111110; B = 8'b10110111; | Outputs: P=%b | Expected: P=%d",
                 1012,
                 
                 P
                 , 
                 
                 11346
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000000; B = 8'b00001101; // Expected: {'P': 2496}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000000; B = 8'b00001101; | Outputs: P=%b | Expected: P=%d",
                 1013,
                 
                 P
                 , 
                 
                 2496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101001; B = 8'b01011001; // Expected: {'P': 20737}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101001; B = 8'b01011001; | Outputs: P=%b | Expected: P=%d",
                 1014,
                 
                 P
                 , 
                 
                 20737
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100001; B = 8'b00111001; // Expected: {'P': 5529}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100001; B = 8'b00111001; | Outputs: P=%b | Expected: P=%d",
                 1015,
                 
                 P
                 , 
                 
                 5529
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001011; B = 8'b01101010; // Expected: {'P': 7950}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001011; B = 8'b01101010; | Outputs: P=%b | Expected: P=%d",
                 1016,
                 
                 P
                 , 
                 
                 7950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001000; B = 8'b10000100; // Expected: {'P': 1056}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001000; B = 8'b10000100; | Outputs: P=%b | Expected: P=%d",
                 1017,
                 
                 P
                 , 
                 
                 1056
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110111; B = 8'b11001001; // Expected: {'P': 49647}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110111; B = 8'b11001001; | Outputs: P=%b | Expected: P=%d",
                 1018,
                 
                 P
                 , 
                 
                 49647
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011101; B = 8'b01000101; // Expected: {'P': 6417}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011101; B = 8'b01000101; | Outputs: P=%b | Expected: P=%d",
                 1019,
                 
                 P
                 , 
                 
                 6417
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111100; B = 8'b10100011; // Expected: {'P': 9780}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111100; B = 8'b10100011; | Outputs: P=%b | Expected: P=%d",
                 1020,
                 
                 P
                 , 
                 
                 9780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100000; B = 8'b11111000; // Expected: {'P': 23808}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100000; B = 8'b11111000; | Outputs: P=%b | Expected: P=%d",
                 1021,
                 
                 P
                 , 
                 
                 23808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111001; B = 8'b10011001; // Expected: {'P': 18513}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111001; B = 8'b10011001; | Outputs: P=%b | Expected: P=%d",
                 1022,
                 
                 P
                 , 
                 
                 18513
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011011; B = 8'b00001011; // Expected: {'P': 1705}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011011; B = 8'b00001011; | Outputs: P=%b | Expected: P=%d",
                 1023,
                 
                 P
                 , 
                 
                 1705
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010010; B = 8'b10110011; // Expected: {'P': 3222}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010010; B = 8'b10110011; | Outputs: P=%b | Expected: P=%d",
                 1024,
                 
                 P
                 , 
                 
                 3222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111000; B = 8'b10110111; // Expected: {'P': 10248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111000; B = 8'b10110111; | Outputs: P=%b | Expected: P=%d",
                 1025,
                 
                 P
                 , 
                 
                 10248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010100; B = 8'b01111000; // Expected: {'P': 2400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010100; B = 8'b01111000; | Outputs: P=%b | Expected: P=%d",
                 1026,
                 
                 P
                 , 
                 
                 2400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000111; B = 8'b01001010; // Expected: {'P': 14726}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000111; B = 8'b01001010; | Outputs: P=%b | Expected: P=%d",
                 1027,
                 
                 P
                 , 
                 
                 14726
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000111; B = 8'b01111101; // Expected: {'P': 24875}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000111; B = 8'b01111101; | Outputs: P=%b | Expected: P=%d",
                 1028,
                 
                 P
                 , 
                 
                 24875
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101110; B = 8'b11110010; // Expected: {'P': 11132}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101110; B = 8'b11110010; | Outputs: P=%b | Expected: P=%d",
                 1029,
                 
                 P
                 , 
                 
                 11132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111111; B = 8'b11001001; // Expected: {'P': 38391}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111111; B = 8'b11001001; | Outputs: P=%b | Expected: P=%d",
                 1030,
                 
                 P
                 , 
                 
                 38391
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100010; B = 8'b01111100; // Expected: {'P': 4216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100010; B = 8'b01111100; | Outputs: P=%b | Expected: P=%d",
                 1031,
                 
                 P
                 , 
                 
                 4216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000110; B = 8'b00111110; // Expected: {'P': 372}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000110; B = 8'b00111110; | Outputs: P=%b | Expected: P=%d",
                 1032,
                 
                 P
                 , 
                 
                 372
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010110; B = 8'b00000101; // Expected: {'P': 750}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010110; B = 8'b00000101; | Outputs: P=%b | Expected: P=%d",
                 1033,
                 
                 P
                 , 
                 
                 750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000011; B = 8'b00010100; // Expected: {'P': 1340}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000011; B = 8'b00010100; | Outputs: P=%b | Expected: P=%d",
                 1034,
                 
                 P
                 , 
                 
                 1340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101110; B = 8'b10100101; // Expected: {'P': 39270}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101110; B = 8'b10100101; | Outputs: P=%b | Expected: P=%d",
                 1035,
                 
                 P
                 , 
                 
                 39270
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010010; B = 8'b11111010; // Expected: {'P': 20500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010010; B = 8'b11111010; | Outputs: P=%b | Expected: P=%d",
                 1036,
                 
                 P
                 , 
                 
                 20500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111111; B = 8'b00100110; // Expected: {'P': 4826}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111111; B = 8'b00100110; | Outputs: P=%b | Expected: P=%d",
                 1037,
                 
                 P
                 , 
                 
                 4826
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111111; B = 8'b01000101; // Expected: {'P': 8763}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111111; B = 8'b01000101; | Outputs: P=%b | Expected: P=%d",
                 1038,
                 
                 P
                 , 
                 
                 8763
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001010; B = 8'b10010011; // Expected: {'P': 29694}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001010; B = 8'b10010011; | Outputs: P=%b | Expected: P=%d",
                 1039,
                 
                 P
                 , 
                 
                 29694
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111110; B = 8'b00000001; // Expected: {'P': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111110; B = 8'b00000001; | Outputs: P=%b | Expected: P=%d",
                 1040,
                 
                 P
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101101; B = 8'b01101011; // Expected: {'P': 18511}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101101; B = 8'b01101011; | Outputs: P=%b | Expected: P=%d",
                 1041,
                 
                 P
                 , 
                 
                 18511
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001001; B = 8'b00000001; // Expected: {'P': 201}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001001; B = 8'b00000001; | Outputs: P=%b | Expected: P=%d",
                 1042,
                 
                 P
                 , 
                 
                 201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000111; B = 8'b01111111; // Expected: {'P': 9017}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000111; B = 8'b01111111; | Outputs: P=%b | Expected: P=%d",
                 1043,
                 
                 P
                 , 
                 
                 9017
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101101; B = 8'b11001000; // Expected: {'P': 47400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101101; B = 8'b11001000; | Outputs: P=%b | Expected: P=%d",
                 1044,
                 
                 P
                 , 
                 
                 47400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011110; B = 8'b01100011; // Expected: {'P': 9306}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011110; B = 8'b01100011; | Outputs: P=%b | Expected: P=%d",
                 1045,
                 
                 P
                 , 
                 
                 9306
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011110; B = 8'b10010111; // Expected: {'P': 4530}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011110; B = 8'b10010111; | Outputs: P=%b | Expected: P=%d",
                 1046,
                 
                 P
                 , 
                 
                 4530
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100001; B = 8'b10010111; // Expected: {'P': 24311}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100001; B = 8'b10010111; | Outputs: P=%b | Expected: P=%d",
                 1047,
                 
                 P
                 , 
                 
                 24311
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110001; B = 8'b00101101; // Expected: {'P': 10845}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110001; B = 8'b00101101; | Outputs: P=%b | Expected: P=%d",
                 1048,
                 
                 P
                 , 
                 
                 10845
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011010; B = 8'b10011100; // Expected: {'P': 4056}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011010; B = 8'b10011100; | Outputs: P=%b | Expected: P=%d",
                 1049,
                 
                 P
                 , 
                 
                 4056
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000001; B = 8'b00100001; // Expected: {'P': 6369}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000001; B = 8'b00100001; | Outputs: P=%b | Expected: P=%d",
                 1050,
                 
                 P
                 , 
                 
                 6369
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111010; B = 8'b01111011; // Expected: {'P': 30750}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111010; B = 8'b01111011; | Outputs: P=%b | Expected: P=%d",
                 1051,
                 
                 P
                 , 
                 
                 30750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110010; B = 8'b01110111; // Expected: {'P': 5950}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110010; B = 8'b01110111; | Outputs: P=%b | Expected: P=%d",
                 1052,
                 
                 P
                 , 
                 
                 5950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011001; B = 8'b11100100; // Expected: {'P': 5700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011001; B = 8'b11100100; | Outputs: P=%b | Expected: P=%d",
                 1053,
                 
                 P
                 , 
                 
                 5700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110100; B = 8'b00010110; // Expected: {'P': 2552}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110100; B = 8'b00010110; | Outputs: P=%b | Expected: P=%d",
                 1054,
                 
                 P
                 , 
                 
                 2552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111001; B = 8'b01111101; // Expected: {'P': 23125}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111001; B = 8'b01111101; | Outputs: P=%b | Expected: P=%d",
                 1055,
                 
                 P
                 , 
                 
                 23125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001101; B = 8'b01000001; // Expected: {'P': 13325}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001101; B = 8'b01000001; | Outputs: P=%b | Expected: P=%d",
                 1056,
                 
                 P
                 , 
                 
                 13325
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101011; B = 8'b00001001; // Expected: {'P': 387}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101011; B = 8'b00001001; | Outputs: P=%b | Expected: P=%d",
                 1057,
                 
                 P
                 , 
                 
                 387
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000101; B = 8'b10000111; // Expected: {'P': 675}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000101; B = 8'b10000111; | Outputs: P=%b | Expected: P=%d",
                 1058,
                 
                 P
                 , 
                 
                 675
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100101; B = 8'b01101101; // Expected: {'P': 24961}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100101; B = 8'b01101101; | Outputs: P=%b | Expected: P=%d",
                 1059,
                 
                 P
                 , 
                 
                 24961
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110110; B = 8'b01110010; // Expected: {'P': 13452}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110110; B = 8'b01110010; | Outputs: P=%b | Expected: P=%d",
                 1060,
                 
                 P
                 , 
                 
                 13452
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100100; B = 8'b11110000; // Expected: {'P': 39360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100100; B = 8'b11110000; | Outputs: P=%b | Expected: P=%d",
                 1061,
                 
                 P
                 , 
                 
                 39360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000110; B = 8'b01101011; // Expected: {'P': 21186}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000110; B = 8'b01101011; | Outputs: P=%b | Expected: P=%d",
                 1062,
                 
                 P
                 , 
                 
                 21186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110000; B = 8'b00010101; // Expected: {'P': 1008}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110000; B = 8'b00010101; | Outputs: P=%b | Expected: P=%d",
                 1063,
                 
                 P
                 , 
                 
                 1008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011111; B = 8'b10110010; // Expected: {'P': 5518}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011111; B = 8'b10110010; | Outputs: P=%b | Expected: P=%d",
                 1064,
                 
                 P
                 , 
                 
                 5518
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001110; B = 8'b10110010; // Expected: {'P': 36668}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001110; B = 8'b10110010; | Outputs: P=%b | Expected: P=%d",
                 1065,
                 
                 P
                 , 
                 
                 36668
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000110; B = 8'b11010000; // Expected: {'P': 14560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000110; B = 8'b11010000; | Outputs: P=%b | Expected: P=%d",
                 1066,
                 
                 P
                 , 
                 
                 14560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100100; B = 8'b11010000; // Expected: {'P': 47424}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100100; B = 8'b11010000; | Outputs: P=%b | Expected: P=%d",
                 1067,
                 
                 P
                 , 
                 
                 47424
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100011; B = 8'b10100111; // Expected: {'P': 16533}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100011; B = 8'b10100111; | Outputs: P=%b | Expected: P=%d",
                 1068,
                 
                 P
                 , 
                 
                 16533
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010101; B = 8'b01110111; // Expected: {'P': 10115}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010101; B = 8'b01110111; | Outputs: P=%b | Expected: P=%d",
                 1069,
                 
                 P
                 , 
                 
                 10115
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100101; B = 8'b10011111; // Expected: {'P': 26235}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100101; B = 8'b10011111; | Outputs: P=%b | Expected: P=%d",
                 1070,
                 
                 P
                 , 
                 
                 26235
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000100; B = 8'b01101000; // Expected: {'P': 13728}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000100; B = 8'b01101000; | Outputs: P=%b | Expected: P=%d",
                 1071,
                 
                 P
                 , 
                 
                 13728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000100; B = 8'b00111000; // Expected: {'P': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000100; B = 8'b00111000; | Outputs: P=%b | Expected: P=%d",
                 1072,
                 
                 P
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000001; B = 8'b11000101; // Expected: {'P': 12805}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000001; B = 8'b11000101; | Outputs: P=%b | Expected: P=%d",
                 1073,
                 
                 P
                 , 
                 
                 12805
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011010; B = 8'b00100010; // Expected: {'P': 5236}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011010; B = 8'b00100010; | Outputs: P=%b | Expected: P=%d",
                 1074,
                 
                 P
                 , 
                 
                 5236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001010; B = 8'b11001100; // Expected: {'P': 15096}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001010; B = 8'b11001100; | Outputs: P=%b | Expected: P=%d",
                 1075,
                 
                 P
                 , 
                 
                 15096
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001010; B = 8'b11111110; // Expected: {'P': 2540}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001010; B = 8'b11111110; | Outputs: P=%b | Expected: P=%d",
                 1076,
                 
                 P
                 , 
                 
                 2540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100100; B = 8'b01010101; // Expected: {'P': 3060}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100100; B = 8'b01010101; | Outputs: P=%b | Expected: P=%d",
                 1077,
                 
                 P
                 , 
                 
                 3060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100001; B = 8'b01101000; // Expected: {'P': 10088}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100001; B = 8'b01101000; | Outputs: P=%b | Expected: P=%d",
                 1078,
                 
                 P
                 , 
                 
                 10088
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001011; B = 8'b11011011; // Expected: {'P': 16425}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001011; B = 8'b11011011; | Outputs: P=%b | Expected: P=%d",
                 1079,
                 
                 P
                 , 
                 
                 16425
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000000; B = 8'b00100110; // Expected: {'P': 2432}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000000; B = 8'b00100110; | Outputs: P=%b | Expected: P=%d",
                 1080,
                 
                 P
                 , 
                 
                 2432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001111; B = 8'b11010100; // Expected: {'P': 43884}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001111; B = 8'b11010100; | Outputs: P=%b | Expected: P=%d",
                 1081,
                 
                 P
                 , 
                 
                 43884
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101011; B = 8'b10000010; // Expected: {'P': 30550}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101011; B = 8'b10000010; | Outputs: P=%b | Expected: P=%d",
                 1082,
                 
                 P
                 , 
                 
                 30550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100110; B = 8'b11110011; // Expected: {'P': 40338}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100110; B = 8'b11110011; | Outputs: P=%b | Expected: P=%d",
                 1083,
                 
                 P
                 , 
                 
                 40338
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010011; B = 8'b11101101; // Expected: {'P': 19671}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010011; B = 8'b11101101; | Outputs: P=%b | Expected: P=%d",
                 1084,
                 
                 P
                 , 
                 
                 19671
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111101; B = 8'b00101111; // Expected: {'P': 11891}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111101; B = 8'b00101111; | Outputs: P=%b | Expected: P=%d",
                 1085,
                 
                 P
                 , 
                 
                 11891
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001101; B = 8'b10100100; // Expected: {'P': 12628}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001101; B = 8'b10100100; | Outputs: P=%b | Expected: P=%d",
                 1086,
                 
                 P
                 , 
                 
                 12628
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010011; B = 8'b00001011; // Expected: {'P': 209}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010011; B = 8'b00001011; | Outputs: P=%b | Expected: P=%d",
                 1087,
                 
                 P
                 , 
                 
                 209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001000; B = 8'b10110011; // Expected: {'P': 24344}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001000; B = 8'b10110011; | Outputs: P=%b | Expected: P=%d",
                 1088,
                 
                 P
                 , 
                 
                 24344
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001000; B = 8'b01101100; // Expected: {'P': 864}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001000; B = 8'b01101100; | Outputs: P=%b | Expected: P=%d",
                 1089,
                 
                 P
                 , 
                 
                 864
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000110; B = 8'b01001111; // Expected: {'P': 10586}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000110; B = 8'b01001111; | Outputs: P=%b | Expected: P=%d",
                 1090,
                 
                 P
                 , 
                 
                 10586
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010110; B = 8'b10000010; // Expected: {'P': 27820}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010110; B = 8'b10000010; | Outputs: P=%b | Expected: P=%d",
                 1091,
                 
                 P
                 , 
                 
                 27820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111001; B = 8'b01100010; // Expected: {'P': 18130}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111001; B = 8'b01100010; | Outputs: P=%b | Expected: P=%d",
                 1092,
                 
                 P
                 , 
                 
                 18130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010011; B = 8'b00011010; // Expected: {'P': 494}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010011; B = 8'b00011010; | Outputs: P=%b | Expected: P=%d",
                 1093,
                 
                 P
                 , 
                 
                 494
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001111; B = 8'b10111111; // Expected: {'P': 2865}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001111; B = 8'b10111111; | Outputs: P=%b | Expected: P=%d",
                 1094,
                 
                 P
                 , 
                 
                 2865
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100001; B = 8'b01010110; // Expected: {'P': 2838}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100001; B = 8'b01010110; | Outputs: P=%b | Expected: P=%d",
                 1095,
                 
                 P
                 , 
                 
                 2838
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100111; B = 8'b10111000; // Expected: {'P': 18952}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100111; B = 8'b10111000; | Outputs: P=%b | Expected: P=%d",
                 1096,
                 
                 P
                 , 
                 
                 18952
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110101; B = 8'b01110001; // Expected: {'P': 20453}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110101; B = 8'b01110001; | Outputs: P=%b | Expected: P=%d",
                 1097,
                 
                 P
                 , 
                 
                 20453
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001010; B = 8'b10001111; // Expected: {'P': 10582}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001010; B = 8'b10001111; | Outputs: P=%b | Expected: P=%d",
                 1098,
                 
                 P
                 , 
                 
                 10582
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100110; B = 8'b01100000; // Expected: {'P': 9792}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100110; B = 8'b01100000; | Outputs: P=%b | Expected: P=%d",
                 1099,
                 
                 P
                 , 
                 
                 9792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000111; B = 8'b00010010; // Expected: {'P': 2430}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000111; B = 8'b00010010; | Outputs: P=%b | Expected: P=%d",
                 1100,
                 
                 P
                 , 
                 
                 2430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110001; B = 8'b10000100; // Expected: {'P': 14916}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110001; B = 8'b10000100; | Outputs: P=%b | Expected: P=%d",
                 1101,
                 
                 P
                 , 
                 
                 14916
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000011; B = 8'b00001011; // Expected: {'P': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000011; B = 8'b00001011; | Outputs: P=%b | Expected: P=%d",
                 1102,
                 
                 P
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101111; B = 8'b01111001; // Expected: {'P': 21175}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101111; B = 8'b01111001; | Outputs: P=%b | Expected: P=%d",
                 1103,
                 
                 P
                 , 
                 
                 21175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001011; B = 8'b01101111; // Expected: {'P': 15429}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001011; B = 8'b01101111; | Outputs: P=%b | Expected: P=%d",
                 1104,
                 
                 P
                 , 
                 
                 15429
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011101; B = 8'b00011111; // Expected: {'P': 4867}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011101; B = 8'b00011111; | Outputs: P=%b | Expected: P=%d",
                 1105,
                 
                 P
                 , 
                 
                 4867
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110111; B = 8'b01011111; // Expected: {'P': 5225}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110111; B = 8'b01011111; | Outputs: P=%b | Expected: P=%d",
                 1106,
                 
                 P
                 , 
                 
                 5225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110011; B = 8'b11111100; // Expected: {'P': 12852}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110011; B = 8'b11111100; | Outputs: P=%b | Expected: P=%d",
                 1107,
                 
                 P
                 , 
                 
                 12852
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100111; B = 8'b00110011; // Expected: {'P': 5253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100111; B = 8'b00110011; | Outputs: P=%b | Expected: P=%d",
                 1108,
                 
                 P
                 , 
                 
                 5253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110000; B = 8'b01000111; // Expected: {'P': 12496}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110000; B = 8'b01000111; | Outputs: P=%b | Expected: P=%d",
                 1109,
                 
                 P
                 , 
                 
                 12496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110100; B = 8'b00010011; // Expected: {'P': 988}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110100; B = 8'b00010011; | Outputs: P=%b | Expected: P=%d",
                 1110,
                 
                 P
                 , 
                 
                 988
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110000; B = 8'b01011000; // Expected: {'P': 9856}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110000; B = 8'b01011000; | Outputs: P=%b | Expected: P=%d",
                 1111,
                 
                 P
                 , 
                 
                 9856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100111; B = 8'b01010001; // Expected: {'P': 8343}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100111; B = 8'b01010001; | Outputs: P=%b | Expected: P=%d",
                 1112,
                 
                 P
                 , 
                 
                 8343
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100110; B = 8'b00000001; // Expected: {'P': 166}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100110; B = 8'b00000001; | Outputs: P=%b | Expected: P=%d",
                 1113,
                 
                 P
                 , 
                 
                 166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010111; B = 8'b01011111; // Expected: {'P': 20425}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010111; B = 8'b01011111; | Outputs: P=%b | Expected: P=%d",
                 1114,
                 
                 P
                 , 
                 
                 20425
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101111; B = 8'b11110001; // Expected: {'P': 26751}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101111; B = 8'b11110001; | Outputs: P=%b | Expected: P=%d",
                 1115,
                 
                 P
                 , 
                 
                 26751
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010100; B = 8'b01101110; // Expected: {'P': 16280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010100; B = 8'b01101110; | Outputs: P=%b | Expected: P=%d",
                 1116,
                 
                 P
                 , 
                 
                 16280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101010; B = 8'b10010100; // Expected: {'P': 6216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101010; B = 8'b10010100; | Outputs: P=%b | Expected: P=%d",
                 1117,
                 
                 P
                 , 
                 
                 6216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010000; B = 8'b11100000; // Expected: {'P': 3584}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010000; B = 8'b11100000; | Outputs: P=%b | Expected: P=%d",
                 1118,
                 
                 P
                 , 
                 
                 3584
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011111; B = 8'b00110100; // Expected: {'P': 11596}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011111; B = 8'b00110100; | Outputs: P=%b | Expected: P=%d",
                 1119,
                 
                 P
                 , 
                 
                 11596
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100001; B = 8'b00011101; // Expected: {'P': 4669}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100001; B = 8'b00011101; | Outputs: P=%b | Expected: P=%d",
                 1120,
                 
                 P
                 , 
                 
                 4669
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111100; B = 8'b01011001; // Expected: {'P': 5340}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111100; B = 8'b01011001; | Outputs: P=%b | Expected: P=%d",
                 1121,
                 
                 P
                 , 
                 
                 5340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010101; B = 8'b01100010; // Expected: {'P': 14602}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010101; B = 8'b01100010; | Outputs: P=%b | Expected: P=%d",
                 1122,
                 
                 P
                 , 
                 
                 14602
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100100; B = 8'b10010010; // Expected: {'P': 5256}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100100; B = 8'b10010010; | Outputs: P=%b | Expected: P=%d",
                 1123,
                 
                 P
                 , 
                 
                 5256
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010111; B = 8'b00111001; // Expected: {'P': 8607}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010111; B = 8'b00111001; | Outputs: P=%b | Expected: P=%d",
                 1124,
                 
                 P
                 , 
                 
                 8607
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010101; B = 8'b11000010; // Expected: {'P': 28906}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010101; B = 8'b11000010; | Outputs: P=%b | Expected: P=%d",
                 1125,
                 
                 P
                 , 
                 
                 28906
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110111; B = 8'b00010000; // Expected: {'P': 2928}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110111; B = 8'b00010000; | Outputs: P=%b | Expected: P=%d",
                 1126,
                 
                 P
                 , 
                 
                 2928
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001100; B = 8'b00011011; // Expected: {'P': 2052}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001100; B = 8'b00011011; | Outputs: P=%b | Expected: P=%d",
                 1127,
                 
                 P
                 , 
                 
                 2052
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101101; B = 8'b10001010; // Expected: {'P': 15042}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101101; B = 8'b10001010; | Outputs: P=%b | Expected: P=%d",
                 1128,
                 
                 P
                 , 
                 
                 15042
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111001; B = 8'b11111111; // Expected: {'P': 14535}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111001; B = 8'b11111111; | Outputs: P=%b | Expected: P=%d",
                 1129,
                 
                 P
                 , 
                 
                 14535
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101100; B = 8'b01100100; // Expected: {'P': 17200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101100; B = 8'b01100100; | Outputs: P=%b | Expected: P=%d",
                 1130,
                 
                 P
                 , 
                 
                 17200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001100; B = 8'b01101101; // Expected: {'P': 15260}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001100; B = 8'b01101101; | Outputs: P=%b | Expected: P=%d",
                 1131,
                 
                 P
                 , 
                 
                 15260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001111; B = 8'b00011000; // Expected: {'P': 3432}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001111; B = 8'b00011000; | Outputs: P=%b | Expected: P=%d",
                 1132,
                 
                 P
                 , 
                 
                 3432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110101; B = 8'b11010011; // Expected: {'P': 11183}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110101; B = 8'b11010011; | Outputs: P=%b | Expected: P=%d",
                 1133,
                 
                 P
                 , 
                 
                 11183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111000; B = 8'b01010100; // Expected: {'P': 10080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111000; B = 8'b01010100; | Outputs: P=%b | Expected: P=%d",
                 1134,
                 
                 P
                 , 
                 
                 10080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000001; B = 8'b10101011; // Expected: {'P': 22059}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000001; B = 8'b10101011; | Outputs: P=%b | Expected: P=%d",
                 1135,
                 
                 P
                 , 
                 
                 22059
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100000; B = 8'b01110111; // Expected: {'P': 19040}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100000; B = 8'b01110111; | Outputs: P=%b | Expected: P=%d",
                 1136,
                 
                 P
                 , 
                 
                 19040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001101; B = 8'b01111011; // Expected: {'P': 25215}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001101; B = 8'b01111011; | Outputs: P=%b | Expected: P=%d",
                 1137,
                 
                 P
                 , 
                 
                 25215
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110010; B = 8'b01001111; // Expected: {'P': 19118}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110010; B = 8'b01001111; | Outputs: P=%b | Expected: P=%d",
                 1138,
                 
                 P
                 , 
                 
                 19118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000111; B = 8'b10011110; // Expected: {'P': 31442}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000111; B = 8'b10011110; | Outputs: P=%b | Expected: P=%d",
                 1139,
                 
                 P
                 , 
                 
                 31442
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110101; B = 8'b00000101; // Expected: {'P': 905}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110101; B = 8'b00000101; | Outputs: P=%b | Expected: P=%d",
                 1140,
                 
                 P
                 , 
                 
                 905
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000010; B = 8'b01001100; // Expected: {'P': 9880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000010; B = 8'b01001100; | Outputs: P=%b | Expected: P=%d",
                 1141,
                 
                 P
                 , 
                 
                 9880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000011; B = 8'b10101001; // Expected: {'P': 11323}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000011; B = 8'b10101001; | Outputs: P=%b | Expected: P=%d",
                 1142,
                 
                 P
                 , 
                 
                 11323
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001001; B = 8'b11001001; // Expected: {'P': 40401}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001001; B = 8'b11001001; | Outputs: P=%b | Expected: P=%d",
                 1143,
                 
                 P
                 , 
                 
                 40401
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101101; B = 8'b11110000; // Expected: {'P': 41520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101101; B = 8'b11110000; | Outputs: P=%b | Expected: P=%d",
                 1144,
                 
                 P
                 , 
                 
                 41520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010010; B = 8'b00001100; // Expected: {'P': 1752}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010010; B = 8'b00001100; | Outputs: P=%b | Expected: P=%d",
                 1145,
                 
                 P
                 , 
                 
                 1752
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001100; B = 8'b00100111; // Expected: {'P': 2964}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001100; B = 8'b00100111; | Outputs: P=%b | Expected: P=%d",
                 1146,
                 
                 P
                 , 
                 
                 2964
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010001; B = 8'b11110000; // Expected: {'P': 50160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010001; B = 8'b11110000; | Outputs: P=%b | Expected: P=%d",
                 1147,
                 
                 P
                 , 
                 
                 50160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011010; B = 8'b11111100; // Expected: {'P': 22680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011010; B = 8'b11111100; | Outputs: P=%b | Expected: P=%d",
                 1148,
                 
                 P
                 , 
                 
                 22680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101001; B = 8'b00000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101001; B = 8'b00000000; | Outputs: P=%b | Expected: P=%d",
                 1149,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111011; B = 8'b00001110; // Expected: {'P': 1722}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111011; B = 8'b00001110; | Outputs: P=%b | Expected: P=%d",
                 1150,
                 
                 P
                 , 
                 
                 1722
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101100; B = 8'b00011010; // Expected: {'P': 2808}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101100; B = 8'b00011010; | Outputs: P=%b | Expected: P=%d",
                 1151,
                 
                 P
                 , 
                 
                 2808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111100; B = 8'b01101100; // Expected: {'P': 13392}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111100; B = 8'b01101100; | Outputs: P=%b | Expected: P=%d",
                 1152,
                 
                 P
                 , 
                 
                 13392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110000; B = 8'b01111100; // Expected: {'P': 29760}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110000; B = 8'b01111100; | Outputs: P=%b | Expected: P=%d",
                 1153,
                 
                 P
                 , 
                 
                 29760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101001; B = 8'b00001101; // Expected: {'P': 3029}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101001; B = 8'b00001101; | Outputs: P=%b | Expected: P=%d",
                 1154,
                 
                 P
                 , 
                 
                 3029
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101111; B = 8'b11010001; // Expected: {'P': 9823}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101111; B = 8'b11010001; | Outputs: P=%b | Expected: P=%d",
                 1155,
                 
                 P
                 , 
                 
                 9823
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010110; B = 8'b10001010; // Expected: {'P': 3036}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010110; B = 8'b10001010; | Outputs: P=%b | Expected: P=%d",
                 1156,
                 
                 P
                 , 
                 
                 3036
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101010; B = 8'b11000001; // Expected: {'P': 32810}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101010; B = 8'b11000001; | Outputs: P=%b | Expected: P=%d",
                 1157,
                 
                 P
                 , 
                 
                 32810
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110011; B = 8'b11010000; // Expected: {'P': 10608}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110011; B = 8'b11010000; | Outputs: P=%b | Expected: P=%d",
                 1158,
                 
                 P
                 , 
                 
                 10608
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100011; B = 8'b11011001; // Expected: {'P': 35371}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100011; B = 8'b11011001; | Outputs: P=%b | Expected: P=%d",
                 1159,
                 
                 P
                 , 
                 
                 35371
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011100; B = 8'b01101101; // Expected: {'P': 17004}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011100; B = 8'b01101101; | Outputs: P=%b | Expected: P=%d",
                 1160,
                 
                 P
                 , 
                 
                 17004
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101000; B = 8'b01101100; // Expected: {'P': 25056}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101000; B = 8'b01101100; | Outputs: P=%b | Expected: P=%d",
                 1161,
                 
                 P
                 , 
                 
                 25056
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011110; B = 8'b10101101; // Expected: {'P': 5190}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011110; B = 8'b10101101; | Outputs: P=%b | Expected: P=%d",
                 1162,
                 
                 P
                 , 
                 
                 5190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001111; B = 8'b11111011; // Expected: {'P': 3765}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001111; B = 8'b11111011; | Outputs: P=%b | Expected: P=%d",
                 1163,
                 
                 P
                 , 
                 
                 3765
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100010; B = 8'b11100001; // Expected: {'P': 50850}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100010; B = 8'b11100001; | Outputs: P=%b | Expected: P=%d",
                 1164,
                 
                 P
                 , 
                 
                 50850
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111011; B = 8'b01010110; // Expected: {'P': 10578}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111011; B = 8'b01010110; | Outputs: P=%b | Expected: P=%d",
                 1165,
                 
                 P
                 , 
                 
                 10578
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011110; B = 8'b10001001; // Expected: {'P': 30414}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011110; B = 8'b10001001; | Outputs: P=%b | Expected: P=%d",
                 1166,
                 
                 P
                 , 
                 
                 30414
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110000; B = 8'b01101000; // Expected: {'P': 11648}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110000; B = 8'b01101000; | Outputs: P=%b | Expected: P=%d",
                 1167,
                 
                 P
                 , 
                 
                 11648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010010; B = 8'b10001101; // Expected: {'P': 2538}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010010; B = 8'b10001101; | Outputs: P=%b | Expected: P=%d",
                 1168,
                 
                 P
                 , 
                 
                 2538
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000001; B = 8'b01010100; // Expected: {'P': 16212}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000001; B = 8'b01010100; | Outputs: P=%b | Expected: P=%d",
                 1169,
                 
                 P
                 , 
                 
                 16212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111111; B = 8'b11000010; // Expected: {'P': 37054}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111111; B = 8'b11000010; | Outputs: P=%b | Expected: P=%d",
                 1170,
                 
                 P
                 , 
                 
                 37054
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100000; B = 8'b00011111; // Expected: {'P': 2976}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100000; B = 8'b00011111; | Outputs: P=%b | Expected: P=%d",
                 1171,
                 
                 P
                 , 
                 
                 2976
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001001; B = 8'b10010100; // Expected: {'P': 10804}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001001; B = 8'b10010100; | Outputs: P=%b | Expected: P=%d",
                 1172,
                 
                 P
                 , 
                 
                 10804
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111111; B = 8'b00111110; // Expected: {'P': 3906}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111111; B = 8'b00111110; | Outputs: P=%b | Expected: P=%d",
                 1173,
                 
                 P
                 , 
                 
                 3906
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101011; B = 8'b01110110; // Expected: {'P': 20178}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101011; B = 8'b01110110; | Outputs: P=%b | Expected: P=%d",
                 1174,
                 
                 P
                 , 
                 
                 20178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110100; B = 8'b10011010; // Expected: {'P': 37576}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110100; B = 8'b10011010; | Outputs: P=%b | Expected: P=%d",
                 1175,
                 
                 P
                 , 
                 
                 37576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100000; B = 8'b01100011; // Expected: {'P': 3168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100000; B = 8'b01100011; | Outputs: P=%b | Expected: P=%d",
                 1176,
                 
                 P
                 , 
                 
                 3168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010100; B = 8'b11111111; // Expected: {'P': 21420}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010100; B = 8'b11111111; | Outputs: P=%b | Expected: P=%d",
                 1177,
                 
                 P
                 , 
                 
                 21420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111101; B = 8'b01011000; // Expected: {'P': 22264}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111101; B = 8'b01011000; | Outputs: P=%b | Expected: P=%d",
                 1178,
                 
                 P
                 , 
                 
                 22264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110111; B = 8'b01111001; // Expected: {'P': 29887}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110111; B = 8'b01111001; | Outputs: P=%b | Expected: P=%d",
                 1179,
                 
                 P
                 , 
                 
                 29887
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001101; B = 8'b00010100; // Expected: {'P': 4100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001101; B = 8'b00010100; | Outputs: P=%b | Expected: P=%d",
                 1180,
                 
                 P
                 , 
                 
                 4100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100000; B = 8'b00110011; // Expected: {'P': 11424}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100000; B = 8'b00110011; | Outputs: P=%b | Expected: P=%d",
                 1181,
                 
                 P
                 , 
                 
                 11424
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101111; B = 8'b10010011; // Expected: {'P': 6909}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101111; B = 8'b10010011; | Outputs: P=%b | Expected: P=%d",
                 1182,
                 
                 P
                 , 
                 
                 6909
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111000; B = 8'b10111101; // Expected: {'P': 22680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111000; B = 8'b10111101; | Outputs: P=%b | Expected: P=%d",
                 1183,
                 
                 P
                 , 
                 
                 22680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011100; B = 8'b01010100; // Expected: {'P': 7728}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011100; B = 8'b01010100; | Outputs: P=%b | Expected: P=%d",
                 1184,
                 
                 P
                 , 
                 
                 7728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111010; B = 8'b11110101; // Expected: {'P': 29890}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111010; B = 8'b11110101; | Outputs: P=%b | Expected: P=%d",
                 1185,
                 
                 P
                 , 
                 
                 29890
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000001; B = 8'b01010100; // Expected: {'P': 10836}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000001; B = 8'b01010100; | Outputs: P=%b | Expected: P=%d",
                 1186,
                 
                 P
                 , 
                 
                 10836
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001110; B = 8'b10110100; // Expected: {'P': 2520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001110; B = 8'b10110100; | Outputs: P=%b | Expected: P=%d",
                 1187,
                 
                 P
                 , 
                 
                 2520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001000; B = 8'b11111000; // Expected: {'P': 17856}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001000; B = 8'b11111000; | Outputs: P=%b | Expected: P=%d",
                 1188,
                 
                 P
                 , 
                 
                 17856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100011; B = 8'b01111101; // Expected: {'P': 12375}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100011; B = 8'b01111101; | Outputs: P=%b | Expected: P=%d",
                 1189,
                 
                 P
                 , 
                 
                 12375
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100100; B = 8'b11010111; // Expected: {'P': 21500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100100; B = 8'b11010111; | Outputs: P=%b | Expected: P=%d",
                 1190,
                 
                 P
                 , 
                 
                 21500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101000; B = 8'b10110000; // Expected: {'P': 7040}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101000; B = 8'b10110000; | Outputs: P=%b | Expected: P=%d",
                 1191,
                 
                 P
                 , 
                 
                 7040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011011; B = 8'b01010110; // Expected: {'P': 13330}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011011; B = 8'b01010110; | Outputs: P=%b | Expected: P=%d",
                 1192,
                 
                 P
                 , 
                 
                 13330
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000010; B = 8'b01010111; // Expected: {'P': 16878}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000010; B = 8'b01010111; | Outputs: P=%b | Expected: P=%d",
                 1193,
                 
                 P
                 , 
                 
                 16878
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010000; B = 8'b01001000; // Expected: {'P': 1152}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010000; B = 8'b01001000; | Outputs: P=%b | Expected: P=%d",
                 1194,
                 
                 P
                 , 
                 
                 1152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100000; B = 8'b10011001; // Expected: {'P': 34272}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100000; B = 8'b10011001; | Outputs: P=%b | Expected: P=%d",
                 1195,
                 
                 P
                 , 
                 
                 34272
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110101; B = 8'b00100010; // Expected: {'P': 6154}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110101; B = 8'b00100010; | Outputs: P=%b | Expected: P=%d",
                 1196,
                 
                 P
                 , 
                 
                 6154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001111; B = 8'b00000001; // Expected: {'P': 143}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001111; B = 8'b00000001; | Outputs: P=%b | Expected: P=%d",
                 1197,
                 
                 P
                 , 
                 
                 143
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011101; B = 8'b11110101; // Expected: {'P': 54145}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011101; B = 8'b11110101; | Outputs: P=%b | Expected: P=%d",
                 1198,
                 
                 P
                 , 
                 
                 54145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010011; B = 8'b10111100; // Expected: {'P': 27636}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010011; B = 8'b10111100; | Outputs: P=%b | Expected: P=%d",
                 1199,
                 
                 P
                 , 
                 
                 27636
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111111; B = 8'b01001101; // Expected: {'P': 19635}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111111; B = 8'b01001101; | Outputs: P=%b | Expected: P=%d",
                 1200,
                 
                 P
                 , 
                 
                 19635
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100000; B = 8'b00010110; // Expected: {'P': 4928}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100000; B = 8'b00010110; | Outputs: P=%b | Expected: P=%d",
                 1201,
                 
                 P
                 , 
                 
                 4928
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010101; B = 8'b10100000; // Expected: {'P': 34080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010101; B = 8'b10100000; | Outputs: P=%b | Expected: P=%d",
                 1202,
                 
                 P
                 , 
                 
                 34080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001011; B = 8'b11001110; // Expected: {'P': 28634}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001011; B = 8'b11001110; | Outputs: P=%b | Expected: P=%d",
                 1203,
                 
                 P
                 , 
                 
                 28634
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100110; B = 8'b01011110; // Expected: {'P': 15604}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100110; B = 8'b01011110; | Outputs: P=%b | Expected: P=%d",
                 1204,
                 
                 P
                 , 
                 
                 15604
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011110; B = 8'b01111011; // Expected: {'P': 3690}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011110; B = 8'b01111011; | Outputs: P=%b | Expected: P=%d",
                 1205,
                 
                 P
                 , 
                 
                 3690
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011001; B = 8'b10000001; // Expected: {'P': 11481}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011001; B = 8'b10000001; | Outputs: P=%b | Expected: P=%d",
                 1206,
                 
                 P
                 , 
                 
                 11481
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010011; B = 8'b11011100; // Expected: {'P': 32340}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010011; B = 8'b11011100; | Outputs: P=%b | Expected: P=%d",
                 1207,
                 
                 P
                 , 
                 
                 32340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011001; B = 8'b11110010; // Expected: {'P': 52514}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011001; B = 8'b11110010; | Outputs: P=%b | Expected: P=%d",
                 1208,
                 
                 P
                 , 
                 
                 52514
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111111; B = 8'b00100110; // Expected: {'P': 7258}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111111; B = 8'b00100110; | Outputs: P=%b | Expected: P=%d",
                 1209,
                 
                 P
                 , 
                 
                 7258
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010001; B = 8'b00000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010001; B = 8'b00000000; | Outputs: P=%b | Expected: P=%d",
                 1210,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111111; B = 8'b00000101; // Expected: {'P': 315}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111111; B = 8'b00000101; | Outputs: P=%b | Expected: P=%d",
                 1211,
                 
                 P
                 , 
                 
                 315
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101011; B = 8'b10110101; // Expected: {'P': 42535}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101011; B = 8'b10110101; | Outputs: P=%b | Expected: P=%d",
                 1212,
                 
                 P
                 , 
                 
                 42535
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001110; B = 8'b01111100; // Expected: {'P': 1736}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001110; B = 8'b01111100; | Outputs: P=%b | Expected: P=%d",
                 1213,
                 
                 P
                 , 
                 
                 1736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101000; B = 8'b11100011; // Expected: {'P': 23608}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101000; B = 8'b11100011; | Outputs: P=%b | Expected: P=%d",
                 1214,
                 
                 P
                 , 
                 
                 23608
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000101; B = 8'b00100110; // Expected: {'P': 2622}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000101; B = 8'b00100110; | Outputs: P=%b | Expected: P=%d",
                 1215,
                 
                 P
                 , 
                 
                 2622
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101101; B = 8'b00001001; // Expected: {'P': 981}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101101; B = 8'b00001001; | Outputs: P=%b | Expected: P=%d",
                 1216,
                 
                 P
                 , 
                 
                 981
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000111; B = 8'b00101110; // Expected: {'P': 9154}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000111; B = 8'b00101110; | Outputs: P=%b | Expected: P=%d",
                 1217,
                 
                 P
                 , 
                 
                 9154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101101; B = 8'b11001100; // Expected: {'P': 22236}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101101; B = 8'b11001100; | Outputs: P=%b | Expected: P=%d",
                 1218,
                 
                 P
                 , 
                 
                 22236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101110; B = 8'b01101110; // Expected: {'P': 5060}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101110; B = 8'b01101110; | Outputs: P=%b | Expected: P=%d",
                 1219,
                 
                 P
                 , 
                 
                 5060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111111; B = 8'b11000100; // Expected: {'P': 24892}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111111; B = 8'b11000100; | Outputs: P=%b | Expected: P=%d",
                 1220,
                 
                 P
                 , 
                 
                 24892
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110111; B = 8'b00100010; // Expected: {'P': 8398}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110111; B = 8'b00100010; | Outputs: P=%b | Expected: P=%d",
                 1221,
                 
                 P
                 , 
                 
                 8398
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001111; B = 8'b11000001; // Expected: {'P': 27599}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001111; B = 8'b11000001; | Outputs: P=%b | Expected: P=%d",
                 1222,
                 
                 P
                 , 
                 
                 27599
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101101; B = 8'b11100100; // Expected: {'P': 54036}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101101; B = 8'b11100100; | Outputs: P=%b | Expected: P=%d",
                 1223,
                 
                 P
                 , 
                 
                 54036
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100001; B = 8'b11111001; // Expected: {'P': 24153}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100001; B = 8'b11111001; | Outputs: P=%b | Expected: P=%d",
                 1224,
                 
                 P
                 , 
                 
                 24153
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110000; B = 8'b01010011; // Expected: {'P': 19920}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110000; B = 8'b01010011; | Outputs: P=%b | Expected: P=%d",
                 1225,
                 
                 P
                 , 
                 
                 19920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001001; B = 8'b00010000; // Expected: {'P': 2192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001001; B = 8'b00010000; | Outputs: P=%b | Expected: P=%d",
                 1226,
                 
                 P
                 , 
                 
                 2192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011101; B = 8'b11101010; // Expected: {'P': 6786}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011101; B = 8'b11101010; | Outputs: P=%b | Expected: P=%d",
                 1227,
                 
                 P
                 , 
                 
                 6786
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000001; B = 8'b01010011; // Expected: {'P': 5395}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000001; B = 8'b01010011; | Outputs: P=%b | Expected: P=%d",
                 1228,
                 
                 P
                 , 
                 
                 5395
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101010; B = 8'b01111101; // Expected: {'P': 29250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101010; B = 8'b01111101; | Outputs: P=%b | Expected: P=%d",
                 1229,
                 
                 P
                 , 
                 
                 29250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001100; B = 8'b11010011; // Expected: {'P': 16036}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001100; B = 8'b11010011; | Outputs: P=%b | Expected: P=%d",
                 1230,
                 
                 P
                 , 
                 
                 16036
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101010; B = 8'b11110111; // Expected: {'P': 10374}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101010; B = 8'b11110111; | Outputs: P=%b | Expected: P=%d",
                 1231,
                 
                 P
                 , 
                 
                 10374
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110110; B = 8'b11100100; // Expected: {'P': 12312}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110110; B = 8'b11100100; | Outputs: P=%b | Expected: P=%d",
                 1232,
                 
                 P
                 , 
                 
                 12312
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100111; B = 8'b11111101; // Expected: {'P': 26059}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100111; B = 8'b11111101; | Outputs: P=%b | Expected: P=%d",
                 1233,
                 
                 P
                 , 
                 
                 26059
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101101; B = 8'b01111110; // Expected: {'P': 21798}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101101; B = 8'b01111110; | Outputs: P=%b | Expected: P=%d",
                 1234,
                 
                 P
                 , 
                 
                 21798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101000; B = 8'b11011110; // Expected: {'P': 8880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101000; B = 8'b11011110; | Outputs: P=%b | Expected: P=%d",
                 1235,
                 
                 P
                 , 
                 
                 8880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110000; B = 8'b01011000; // Expected: {'P': 4224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110000; B = 8'b01011000; | Outputs: P=%b | Expected: P=%d",
                 1236,
                 
                 P
                 , 
                 
                 4224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111001; B = 8'b10000100; // Expected: {'P': 7524}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111001; B = 8'b10000100; | Outputs: P=%b | Expected: P=%d",
                 1237,
                 
                 P
                 , 
                 
                 7524
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001110; B = 8'b00101000; // Expected: {'P': 5680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001110; B = 8'b00101000; | Outputs: P=%b | Expected: P=%d",
                 1238,
                 
                 P
                 , 
                 
                 5680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111010; B = 8'b11011111; // Expected: {'P': 41478}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111010; B = 8'b11011111; | Outputs: P=%b | Expected: P=%d",
                 1239,
                 
                 P
                 , 
                 
                 41478
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001110; B = 8'b11100010; // Expected: {'P': 17628}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001110; B = 8'b11100010; | Outputs: P=%b | Expected: P=%d",
                 1240,
                 
                 P
                 , 
                 
                 17628
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101000; B = 8'b00111110; // Expected: {'P': 2480}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101000; B = 8'b00111110; | Outputs: P=%b | Expected: P=%d",
                 1241,
                 
                 P
                 , 
                 
                 2480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101001; B = 8'b11101111; // Expected: {'P': 55687}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101001; B = 8'b11101111; | Outputs: P=%b | Expected: P=%d",
                 1242,
                 
                 P
                 , 
                 
                 55687
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000010; B = 8'b01111101; // Expected: {'P': 8250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000010; B = 8'b01111101; | Outputs: P=%b | Expected: P=%d",
                 1243,
                 
                 P
                 , 
                 
                 8250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111101; B = 8'b11011000; // Expected: {'P': 40824}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111101; B = 8'b11011000; | Outputs: P=%b | Expected: P=%d",
                 1244,
                 
                 P
                 , 
                 
                 40824
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000011; B = 8'b10110000; // Expected: {'P': 34320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000011; B = 8'b10110000; | Outputs: P=%b | Expected: P=%d",
                 1245,
                 
                 P
                 , 
                 
                 34320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000011; B = 8'b11001000; // Expected: {'P': 39000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000011; B = 8'b11001000; | Outputs: P=%b | Expected: P=%d",
                 1246,
                 
                 P
                 , 
                 
                 39000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000001; B = 8'b11010110; // Expected: {'P': 41302}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000001; B = 8'b11010110; | Outputs: P=%b | Expected: P=%d",
                 1247,
                 
                 P
                 , 
                 
                 41302
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001001; B = 8'b01110000; // Expected: {'P': 8176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001001; B = 8'b01110000; | Outputs: P=%b | Expected: P=%d",
                 1248,
                 
                 P
                 , 
                 
                 8176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001011; B = 8'b01001010; // Expected: {'P': 15022}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001011; B = 8'b01001010; | Outputs: P=%b | Expected: P=%d",
                 1249,
                 
                 P
                 , 
                 
                 15022
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111111; B = 8'b00100010; // Expected: {'P': 6494}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111111; B = 8'b00100010; | Outputs: P=%b | Expected: P=%d",
                 1250,
                 
                 P
                 , 
                 
                 6494
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100110; B = 8'b11101010; // Expected: {'P': 8892}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100110; B = 8'b11101010; | Outputs: P=%b | Expected: P=%d",
                 1251,
                 
                 P
                 , 
                 
                 8892
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000110; B = 8'b00111000; // Expected: {'P': 7504}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000110; B = 8'b00111000; | Outputs: P=%b | Expected: P=%d",
                 1252,
                 
                 P
                 , 
                 
                 7504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010010; B = 8'b10001011; // Expected: {'P': 11398}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010010; B = 8'b10001011; | Outputs: P=%b | Expected: P=%d",
                 1253,
                 
                 P
                 , 
                 
                 11398
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110110; B = 8'b10101001; // Expected: {'P': 30758}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110110; B = 8'b10101001; | Outputs: P=%b | Expected: P=%d",
                 1254,
                 
                 P
                 , 
                 
                 30758
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011111; B = 8'b00011001; // Expected: {'P': 5575}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011111; B = 8'b00011001; | Outputs: P=%b | Expected: P=%d",
                 1255,
                 
                 P
                 , 
                 
                 5575
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000101; B = 8'b01110000; // Expected: {'P': 14896}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000101; B = 8'b01110000; | Outputs: P=%b | Expected: P=%d",
                 1256,
                 
                 P
                 , 
                 
                 14896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111011; B = 8'b11110111; // Expected: {'P': 61997}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111011; B = 8'b11110111; | Outputs: P=%b | Expected: P=%d",
                 1257,
                 
                 P
                 , 
                 
                 61997
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100111; B = 8'b01000000; // Expected: {'P': 6592}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100111; B = 8'b01000000; | Outputs: P=%b | Expected: P=%d",
                 1258,
                 
                 P
                 , 
                 
                 6592
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101101; B = 8'b00011010; // Expected: {'P': 6162}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101101; B = 8'b00011010; | Outputs: P=%b | Expected: P=%d",
                 1259,
                 
                 P
                 , 
                 
                 6162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101111; B = 8'b00011010; // Expected: {'P': 1222}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101111; B = 8'b00011010; | Outputs: P=%b | Expected: P=%d",
                 1260,
                 
                 P
                 , 
                 
                 1222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000110; B = 8'b01110111; // Expected: {'P': 23562}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000110; B = 8'b01110111; | Outputs: P=%b | Expected: P=%d",
                 1261,
                 
                 P
                 , 
                 
                 23562
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101100; B = 8'b11001000; // Expected: {'P': 8800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101100; B = 8'b11001000; | Outputs: P=%b | Expected: P=%d",
                 1262,
                 
                 P
                 , 
                 
                 8800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111111; B = 8'b10111111; // Expected: {'P': 12033}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111111; B = 8'b10111111; | Outputs: P=%b | Expected: P=%d",
                 1263,
                 
                 P
                 , 
                 
                 12033
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110010; B = 8'b10111000; // Expected: {'P': 44528}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110010; B = 8'b10111000; | Outputs: P=%b | Expected: P=%d",
                 1264,
                 
                 P
                 , 
                 
                 44528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111101; B = 8'b00001000; // Expected: {'P': 2024}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111101; B = 8'b00001000; | Outputs: P=%b | Expected: P=%d",
                 1265,
                 
                 P
                 , 
                 
                 2024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010111; B = 8'b01010001; // Expected: {'P': 1863}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010111; B = 8'b01010001; | Outputs: P=%b | Expected: P=%d",
                 1266,
                 
                 P
                 , 
                 
                 1863
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011001; B = 8'b10110111; // Expected: {'P': 27999}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011001; B = 8'b10110111; | Outputs: P=%b | Expected: P=%d",
                 1267,
                 
                 P
                 , 
                 
                 27999
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110100; B = 8'b10100000; // Expected: {'P': 28800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110100; B = 8'b10100000; | Outputs: P=%b | Expected: P=%d",
                 1268,
                 
                 P
                 , 
                 
                 28800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000010; B = 8'b11011111; // Expected: {'P': 14718}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000010; B = 8'b11011111; | Outputs: P=%b | Expected: P=%d",
                 1269,
                 
                 P
                 , 
                 
                 14718
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010011; B = 8'b10010100; // Expected: {'P': 12284}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010011; B = 8'b10010100; | Outputs: P=%b | Expected: P=%d",
                 1270,
                 
                 P
                 , 
                 
                 12284
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000001; B = 8'b01000000; // Expected: {'P': 12352}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000001; B = 8'b01000000; | Outputs: P=%b | Expected: P=%d",
                 1271,
                 
                 P
                 , 
                 
                 12352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111001; B = 8'b10110100; // Expected: {'P': 33300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111001; B = 8'b10110100; | Outputs: P=%b | Expected: P=%d",
                 1272,
                 
                 P
                 , 
                 
                 33300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110110; B = 8'b00010101; // Expected: {'P': 5166}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110110; B = 8'b00010101; | Outputs: P=%b | Expected: P=%d",
                 1273,
                 
                 P
                 , 
                 
                 5166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111100; B = 8'b01000100; // Expected: {'P': 8432}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111100; B = 8'b01000100; | Outputs: P=%b | Expected: P=%d",
                 1274,
                 
                 P
                 , 
                 
                 8432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011111; B = 8'b00111001; // Expected: {'P': 9063}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011111; B = 8'b00111001; | Outputs: P=%b | Expected: P=%d",
                 1275,
                 
                 P
                 , 
                 
                 9063
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000100; B = 8'b11000001; // Expected: {'P': 25476}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000100; B = 8'b11000001; | Outputs: P=%b | Expected: P=%d",
                 1276,
                 
                 P
                 , 
                 
                 25476
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101111; B = 8'b10010100; // Expected: {'P': 6956}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101111; B = 8'b10010100; | Outputs: P=%b | Expected: P=%d",
                 1277,
                 
                 P
                 , 
                 
                 6956
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000010; B = 8'b11010001; // Expected: {'P': 40546}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000010; B = 8'b11010001; | Outputs: P=%b | Expected: P=%d",
                 1278,
                 
                 P
                 , 
                 
                 40546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100011; B = 8'b11011010; // Expected: {'P': 21582}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100011; B = 8'b11011010; | Outputs: P=%b | Expected: P=%d",
                 1279,
                 
                 P
                 , 
                 
                 21582
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101110; B = 8'b00000010; // Expected: {'P': 220}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101110; B = 8'b00000010; | Outputs: P=%b | Expected: P=%d",
                 1280,
                 
                 P
                 , 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110000; B = 8'b10011011; // Expected: {'P': 27280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110000; B = 8'b10011011; | Outputs: P=%b | Expected: P=%d",
                 1281,
                 
                 P
                 , 
                 
                 27280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010110; B = 8'b00111101; // Expected: {'P': 5246}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010110; B = 8'b00111101; | Outputs: P=%b | Expected: P=%d",
                 1282,
                 
                 P
                 , 
                 
                 5246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110100; B = 8'b00101000; // Expected: {'P': 2080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110100; B = 8'b00101000; | Outputs: P=%b | Expected: P=%d",
                 1283,
                 
                 P
                 , 
                 
                 2080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111001; B = 8'b00101101; // Expected: {'P': 2565}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111001; B = 8'b00101101; | Outputs: P=%b | Expected: P=%d",
                 1284,
                 
                 P
                 , 
                 
                 2565
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010001; B = 8'b11101000; // Expected: {'P': 48488}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010001; B = 8'b11101000; | Outputs: P=%b | Expected: P=%d",
                 1285,
                 
                 P
                 , 
                 
                 48488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110110; B = 8'b10010011; // Expected: {'P': 7938}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110110; B = 8'b10010011; | Outputs: P=%b | Expected: P=%d",
                 1286,
                 
                 P
                 , 
                 
                 7938
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101010; B = 8'b10100110; // Expected: {'P': 17596}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101010; B = 8'b10100110; | Outputs: P=%b | Expected: P=%d",
                 1287,
                 
                 P
                 , 
                 
                 17596
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010001; B = 8'b01101000; // Expected: {'P': 8424}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010001; B = 8'b01101000; | Outputs: P=%b | Expected: P=%d",
                 1288,
                 
                 P
                 , 
                 
                 8424
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110100; B = 8'b00001000; // Expected: {'P': 1440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110100; B = 8'b00001000; | Outputs: P=%b | Expected: P=%d",
                 1289,
                 
                 P
                 , 
                 
                 1440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101010; B = 8'b00101001; // Expected: {'P': 4346}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101010; B = 8'b00101001; | Outputs: P=%b | Expected: P=%d",
                 1290,
                 
                 P
                 , 
                 
                 4346
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100001; B = 8'b00011010; // Expected: {'P': 858}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100001; B = 8'b00011010; | Outputs: P=%b | Expected: P=%d",
                 1291,
                 
                 P
                 , 
                 
                 858
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100111; B = 8'b10111001; // Expected: {'P': 30895}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100111; B = 8'b10111001; | Outputs: P=%b | Expected: P=%d",
                 1292,
                 
                 P
                 , 
                 
                 30895
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100011; B = 8'b01000101; // Expected: {'P': 15663}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100011; B = 8'b01000101; | Outputs: P=%b | Expected: P=%d",
                 1293,
                 
                 P
                 , 
                 
                 15663
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100101; B = 8'b00010001; // Expected: {'P': 629}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100101; B = 8'b00010001; | Outputs: P=%b | Expected: P=%d",
                 1294,
                 
                 P
                 , 
                 
                 629
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110101; B = 8'b01101000; // Expected: {'P': 25480}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110101; B = 8'b01101000; | Outputs: P=%b | Expected: P=%d",
                 1295,
                 
                 P
                 , 
                 
                 25480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011001; B = 8'b01001000; // Expected: {'P': 11016}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011001; B = 8'b01001000; | Outputs: P=%b | Expected: P=%d",
                 1296,
                 
                 P
                 , 
                 
                 11016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001110; B = 8'b01101011; // Expected: {'P': 22042}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001110; B = 8'b01101011; | Outputs: P=%b | Expected: P=%d",
                 1297,
                 
                 P
                 , 
                 
                 22042
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001101; B = 8'b01001000; // Expected: {'P': 10152}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001101; B = 8'b01001000; | Outputs: P=%b | Expected: P=%d",
                 1298,
                 
                 P
                 , 
                 
                 10152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100010; B = 8'b11001000; // Expected: {'P': 19600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100010; B = 8'b11001000; | Outputs: P=%b | Expected: P=%d",
                 1299,
                 
                 P
                 , 
                 
                 19600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000100; B = 8'b10011110; // Expected: {'P': 10744}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000100; B = 8'b10011110; | Outputs: P=%b | Expected: P=%d",
                 1300,
                 
                 P
                 , 
                 
                 10744
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100011; B = 8'b11001110; // Expected: {'P': 46762}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100011; B = 8'b11001110; | Outputs: P=%b | Expected: P=%d",
                 1301,
                 
                 P
                 , 
                 
                 46762
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011001; B = 8'b00010110; // Expected: {'P': 4774}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011001; B = 8'b00010110; | Outputs: P=%b | Expected: P=%d",
                 1302,
                 
                 P
                 , 
                 
                 4774
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010010; B = 8'b10000011; // Expected: {'P': 19126}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010010; B = 8'b10000011; | Outputs: P=%b | Expected: P=%d",
                 1303,
                 
                 P
                 , 
                 
                 19126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010000; B = 8'b10111000; // Expected: {'P': 14720}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010000; B = 8'b10111000; | Outputs: P=%b | Expected: P=%d",
                 1304,
                 
                 P
                 , 
                 
                 14720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001101; B = 8'b00010011; // Expected: {'P': 247}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001101; B = 8'b00010011; | Outputs: P=%b | Expected: P=%d",
                 1305,
                 
                 P
                 , 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011001; B = 8'b00011101; // Expected: {'P': 6293}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011001; B = 8'b00011101; | Outputs: P=%b | Expected: P=%d",
                 1306,
                 
                 P
                 , 
                 
                 6293
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000000; B = 8'b10101010; // Expected: {'P': 10880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000000; B = 8'b10101010; | Outputs: P=%b | Expected: P=%d",
                 1307,
                 
                 P
                 , 
                 
                 10880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111100; B = 8'b01101010; // Expected: {'P': 26712}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111100; B = 8'b01101010; | Outputs: P=%b | Expected: P=%d",
                 1308,
                 
                 P
                 , 
                 
                 26712
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000100; B = 8'b10111111; // Expected: {'P': 12988}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000100; B = 8'b10111111; | Outputs: P=%b | Expected: P=%d",
                 1309,
                 
                 P
                 , 
                 
                 12988
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100010; B = 8'b10110011; // Expected: {'P': 17542}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100010; B = 8'b10110011; | Outputs: P=%b | Expected: P=%d",
                 1310,
                 
                 P
                 , 
                 
                 17542
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010100; B = 8'b10110001; // Expected: {'P': 26196}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010100; B = 8'b10110001; | Outputs: P=%b | Expected: P=%d",
                 1311,
                 
                 P
                 , 
                 
                 26196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001100; B = 8'b11001100; // Expected: {'P': 28560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001100; B = 8'b11001100; | Outputs: P=%b | Expected: P=%d",
                 1312,
                 
                 P
                 , 
                 
                 28560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100100; B = 8'b11011111; // Expected: {'P': 50844}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100100; B = 8'b11011111; | Outputs: P=%b | Expected: P=%d",
                 1313,
                 
                 P
                 , 
                 
                 50844
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100101; B = 8'b00010001; // Expected: {'P': 2805}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100101; B = 8'b00010001; | Outputs: P=%b | Expected: P=%d",
                 1314,
                 
                 P
                 , 
                 
                 2805
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001001; B = 8'b01000100; // Expected: {'P': 4964}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001001; B = 8'b01000100; | Outputs: P=%b | Expected: P=%d",
                 1315,
                 
                 P
                 , 
                 
                 4964
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001001; B = 8'b10011101; // Expected: {'P': 21509}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001001; B = 8'b10011101; | Outputs: P=%b | Expected: P=%d",
                 1316,
                 
                 P
                 , 
                 
                 21509
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101110; B = 8'b10011101; // Expected: {'P': 17270}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101110; B = 8'b10011101; | Outputs: P=%b | Expected: P=%d",
                 1317,
                 
                 P
                 , 
                 
                 17270
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110010; B = 8'b01001100; // Expected: {'P': 13528}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110010; B = 8'b01001100; | Outputs: P=%b | Expected: P=%d",
                 1318,
                 
                 P
                 , 
                 
                 13528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010101; B = 8'b10011010; // Expected: {'P': 22946}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010101; B = 8'b10011010; | Outputs: P=%b | Expected: P=%d",
                 1319,
                 
                 P
                 , 
                 
                 22946
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111110; B = 8'b00111110; // Expected: {'P': 11780}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111110; B = 8'b00111110; | Outputs: P=%b | Expected: P=%d",
                 1320,
                 
                 P
                 , 
                 
                 11780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011011; B = 8'b01101100; // Expected: {'P': 9828}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011011; B = 8'b01101100; | Outputs: P=%b | Expected: P=%d",
                 1321,
                 
                 P
                 , 
                 
                 9828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111100; B = 8'b11111010; // Expected: {'P': 31000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111100; B = 8'b11111010; | Outputs: P=%b | Expected: P=%d",
                 1322,
                 
                 P
                 , 
                 
                 31000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101001; B = 8'b10110101; // Expected: {'P': 19005}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101001; B = 8'b10110101; | Outputs: P=%b | Expected: P=%d",
                 1323,
                 
                 P
                 , 
                 
                 19005
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101110; B = 8'b01110111; // Expected: {'P': 5474}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101110; B = 8'b01110111; | Outputs: P=%b | Expected: P=%d",
                 1324,
                 
                 P
                 , 
                 
                 5474
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101010; B = 8'b01111101; // Expected: {'P': 5250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101010; B = 8'b01111101; | Outputs: P=%b | Expected: P=%d",
                 1325,
                 
                 P
                 , 
                 
                 5250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111000; B = 8'b10000101; // Expected: {'P': 24472}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111000; B = 8'b10000101; | Outputs: P=%b | Expected: P=%d",
                 1326,
                 
                 P
                 , 
                 
                 24472
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101011; B = 8'b11111110; // Expected: {'P': 10922}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101011; B = 8'b11111110; | Outputs: P=%b | Expected: P=%d",
                 1327,
                 
                 P
                 , 
                 
                 10922
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011011; B = 8'b10110000; // Expected: {'P': 38544}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011011; B = 8'b10110000; | Outputs: P=%b | Expected: P=%d",
                 1328,
                 
                 P
                 , 
                 
                 38544
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110101; B = 8'b11001111; // Expected: {'P': 24219}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110101; B = 8'b11001111; | Outputs: P=%b | Expected: P=%d",
                 1329,
                 
                 P
                 , 
                 
                 24219
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011000; B = 8'b11111110; // Expected: {'P': 6096}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011000; B = 8'b11111110; | Outputs: P=%b | Expected: P=%d",
                 1330,
                 
                 P
                 , 
                 
                 6096
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110010; B = 8'b10010100; // Expected: {'P': 16872}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110010; B = 8'b10010100; | Outputs: P=%b | Expected: P=%d",
                 1331,
                 
                 P
                 , 
                 
                 16872
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110111; B = 8'b01100100; // Expected: {'P': 11900}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110111; B = 8'b01100100; | Outputs: P=%b | Expected: P=%d",
                 1332,
                 
                 P
                 , 
                 
                 11900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001000; B = 8'b01011100; // Expected: {'P': 6624}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001000; B = 8'b01011100; | Outputs: P=%b | Expected: P=%d",
                 1333,
                 
                 P
                 , 
                 
                 6624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101001; B = 8'b10110011; // Expected: {'P': 30251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101001; B = 8'b10110011; | Outputs: P=%b | Expected: P=%d",
                 1334,
                 
                 P
                 , 
                 
                 30251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100000; B = 8'b11111000; // Expected: {'P': 39680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100000; B = 8'b11111000; | Outputs: P=%b | Expected: P=%d",
                 1335,
                 
                 P
                 , 
                 
                 39680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000001; B = 8'b00110101; // Expected: {'P': 10229}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000001; B = 8'b00110101; | Outputs: P=%b | Expected: P=%d",
                 1336,
                 
                 P
                 , 
                 
                 10229
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111011; B = 8'b00010001; // Expected: {'P': 2091}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111011; B = 8'b00010001; | Outputs: P=%b | Expected: P=%d",
                 1337,
                 
                 P
                 , 
                 
                 2091
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110011; B = 8'b10110011; // Expected: {'P': 9129}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110011; B = 8'b10110011; | Outputs: P=%b | Expected: P=%d",
                 1338,
                 
                 P
                 , 
                 
                 9129
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100111; B = 8'b11101011; // Expected: {'P': 39245}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100111; B = 8'b11101011; | Outputs: P=%b | Expected: P=%d",
                 1339,
                 
                 P
                 , 
                 
                 39245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001100; B = 8'b01101111; // Expected: {'P': 22644}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001100; B = 8'b01101111; | Outputs: P=%b | Expected: P=%d",
                 1340,
                 
                 P
                 , 
                 
                 22644
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101110; B = 8'b01001101; // Expected: {'P': 8470}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101110; B = 8'b01001101; | Outputs: P=%b | Expected: P=%d",
                 1341,
                 
                 P
                 , 
                 
                 8470
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111100; B = 8'b10110001; // Expected: {'P': 44604}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111100; B = 8'b10110001; | Outputs: P=%b | Expected: P=%d",
                 1342,
                 
                 P
                 , 
                 
                 44604
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000000; B = 8'b01100101; // Expected: {'P': 19392}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000000; B = 8'b01100101; | Outputs: P=%b | Expected: P=%d",
                 1343,
                 
                 P
                 , 
                 
                 19392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010011; B = 8'b00111100; // Expected: {'P': 8820}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010011; B = 8'b00111100; | Outputs: P=%b | Expected: P=%d",
                 1344,
                 
                 P
                 , 
                 
                 8820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000010; B = 8'b10101101; // Expected: {'P': 33562}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000010; B = 8'b10101101; | Outputs: P=%b | Expected: P=%d",
                 1345,
                 
                 P
                 , 
                 
                 33562
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110100; B = 8'b10110011; // Expected: {'P': 43676}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110100; B = 8'b10110011; | Outputs: P=%b | Expected: P=%d",
                 1346,
                 
                 P
                 , 
                 
                 43676
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001101; B = 8'b11100010; // Expected: {'P': 17402}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001101; B = 8'b11100010; | Outputs: P=%b | Expected: P=%d",
                 1347,
                 
                 P
                 , 
                 
                 17402
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011100; B = 8'b00001111; // Expected: {'P': 420}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011100; B = 8'b00001111; | Outputs: P=%b | Expected: P=%d",
                 1348,
                 
                 P
                 , 
                 
                 420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010011; B = 8'b01010100; // Expected: {'P': 1596}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010011; B = 8'b01010100; | Outputs: P=%b | Expected: P=%d",
                 1349,
                 
                 P
                 , 
                 
                 1596
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110111; B = 8'b00111000; // Expected: {'P': 6664}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110111; B = 8'b00111000; | Outputs: P=%b | Expected: P=%d",
                 1350,
                 
                 P
                 , 
                 
                 6664
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000001; B = 8'b11101111; // Expected: {'P': 46127}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000001; B = 8'b11101111; | Outputs: P=%b | Expected: P=%d",
                 1351,
                 
                 P
                 , 
                 
                 46127
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100111; B = 8'b01101110; // Expected: {'P': 11330}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100111; B = 8'b01101110; | Outputs: P=%b | Expected: P=%d",
                 1352,
                 
                 P
                 , 
                 
                 11330
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010101; B = 8'b10010101; // Expected: {'P': 12665}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010101; B = 8'b10010101; | Outputs: P=%b | Expected: P=%d",
                 1353,
                 
                 P
                 , 
                 
                 12665
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100011; B = 8'b11011000; // Expected: {'P': 35208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100011; B = 8'b11011000; | Outputs: P=%b | Expected: P=%d",
                 1354,
                 
                 P
                 , 
                 
                 35208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111001; B = 8'b00000110; // Expected: {'P': 726}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111001; B = 8'b00000110; | Outputs: P=%b | Expected: P=%d",
                 1355,
                 
                 P
                 , 
                 
                 726
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100000; B = 8'b01011010; // Expected: {'P': 14400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100000; B = 8'b01011010; | Outputs: P=%b | Expected: P=%d",
                 1356,
                 
                 P
                 , 
                 
                 14400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111101; B = 8'b10100010; // Expected: {'P': 9882}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111101; B = 8'b10100010; | Outputs: P=%b | Expected: P=%d",
                 1357,
                 
                 P
                 , 
                 
                 9882
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010110; B = 8'b10010011; // Expected: {'P': 12642}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010110; B = 8'b10010011; | Outputs: P=%b | Expected: P=%d",
                 1358,
                 
                 P
                 , 
                 
                 12642
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111100; B = 8'b11011100; // Expected: {'P': 13200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111100; B = 8'b11011100; | Outputs: P=%b | Expected: P=%d",
                 1359,
                 
                 P
                 , 
                 
                 13200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100000; B = 8'b10001001; // Expected: {'P': 4384}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100000; B = 8'b10001001; | Outputs: P=%b | Expected: P=%d",
                 1360,
                 
                 P
                 , 
                 
                 4384
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111110; B = 8'b01111011; // Expected: {'P': 23370}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111110; B = 8'b01111011; | Outputs: P=%b | Expected: P=%d",
                 1361,
                 
                 P
                 , 
                 
                 23370
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000101; B = 8'b11100000; // Expected: {'P': 1120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000101; B = 8'b11100000; | Outputs: P=%b | Expected: P=%d",
                 1362,
                 
                 P
                 , 
                 
                 1120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111011; B = 8'b00001101; // Expected: {'P': 767}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111011; B = 8'b00001101; | Outputs: P=%b | Expected: P=%d",
                 1363,
                 
                 P
                 , 
                 
                 767
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100110; B = 8'b11111101; // Expected: {'P': 41998}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100110; B = 8'b11111101; | Outputs: P=%b | Expected: P=%d",
                 1364,
                 
                 P
                 , 
                 
                 41998
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000010; B = 8'b10110011; // Expected: {'P': 11814}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000010; B = 8'b10110011; | Outputs: P=%b | Expected: P=%d",
                 1365,
                 
                 P
                 , 
                 
                 11814
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011101; B = 8'b00000010; // Expected: {'P': 186}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011101; B = 8'b00000010; | Outputs: P=%b | Expected: P=%d",
                 1366,
                 
                 P
                 , 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001000; B = 8'b01010011; // Expected: {'P': 664}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001000; B = 8'b01010011; | Outputs: P=%b | Expected: P=%d",
                 1367,
                 
                 P
                 , 
                 
                 664
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111000; B = 8'b11011000; // Expected: {'P': 39744}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111000; B = 8'b11011000; | Outputs: P=%b | Expected: P=%d",
                 1368,
                 
                 P
                 , 
                 
                 39744
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001111; B = 8'b11101111; // Expected: {'P': 49473}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001111; B = 8'b11101111; | Outputs: P=%b | Expected: P=%d",
                 1369,
                 
                 P
                 , 
                 
                 49473
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111101; B = 8'b00101001; // Expected: {'P': 7749}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111101; B = 8'b00101001; | Outputs: P=%b | Expected: P=%d",
                 1370,
                 
                 P
                 , 
                 
                 7749
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010110; B = 8'b10110000; // Expected: {'P': 37664}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010110; B = 8'b10110000; | Outputs: P=%b | Expected: P=%d",
                 1371,
                 
                 P
                 , 
                 
                 37664
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011010; B = 8'b00001010; // Expected: {'P': 2180}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011010; B = 8'b00001010; | Outputs: P=%b | Expected: P=%d",
                 1372,
                 
                 P
                 , 
                 
                 2180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001001; B = 8'b11000010; // Expected: {'P': 1746}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001001; B = 8'b11000010; | Outputs: P=%b | Expected: P=%d",
                 1373,
                 
                 P
                 , 
                 
                 1746
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010100; B = 8'b00001110; // Expected: {'P': 1176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010100; B = 8'b00001110; | Outputs: P=%b | Expected: P=%d",
                 1374,
                 
                 P
                 , 
                 
                 1176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010011; B = 8'b00110101; // Expected: {'P': 4399}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010011; B = 8'b00110101; | Outputs: P=%b | Expected: P=%d",
                 1375,
                 
                 P
                 , 
                 
                 4399
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001111; B = 8'b01111011; // Expected: {'P': 25461}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001111; B = 8'b01111011; | Outputs: P=%b | Expected: P=%d",
                 1376,
                 
                 P
                 , 
                 
                 25461
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111110; B = 8'b10111010; // Expected: {'P': 47244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111110; B = 8'b10111010; | Outputs: P=%b | Expected: P=%d",
                 1377,
                 
                 P
                 , 
                 
                 47244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011011; B = 8'b01001000; // Expected: {'P': 1944}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011011; B = 8'b01001000; | Outputs: P=%b | Expected: P=%d",
                 1378,
                 
                 P
                 , 
                 
                 1944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110010; B = 8'b01101001; // Expected: {'P': 5250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110010; B = 8'b01101001; | Outputs: P=%b | Expected: P=%d",
                 1379,
                 
                 P
                 , 
                 
                 5250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011100; B = 8'b00001000; // Expected: {'P': 1760}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011100; B = 8'b00001000; | Outputs: P=%b | Expected: P=%d",
                 1380,
                 
                 P
                 , 
                 
                 1760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011100; B = 8'b11101110; // Expected: {'P': 21896}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011100; B = 8'b11101110; | Outputs: P=%b | Expected: P=%d",
                 1381,
                 
                 P
                 , 
                 
                 21896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010001; B = 8'b00110101; // Expected: {'P': 11077}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010001; B = 8'b00110101; | Outputs: P=%b | Expected: P=%d",
                 1382,
                 
                 P
                 , 
                 
                 11077
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010101; B = 8'b01001001; // Expected: {'P': 1533}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010101; B = 8'b01001001; | Outputs: P=%b | Expected: P=%d",
                 1383,
                 
                 P
                 , 
                 
                 1533
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111010; B = 8'b00101101; // Expected: {'P': 2610}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111010; B = 8'b00101101; | Outputs: P=%b | Expected: P=%d",
                 1384,
                 
                 P
                 , 
                 
                 2610
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111110; B = 8'b10001000; // Expected: {'P': 17136}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111110; B = 8'b10001000; | Outputs: P=%b | Expected: P=%d",
                 1385,
                 
                 P
                 , 
                 
                 17136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110010; B = 8'b00000011; // Expected: {'P': 150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110010; B = 8'b00000011; | Outputs: P=%b | Expected: P=%d",
                 1386,
                 
                 P
                 , 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000111; B = 8'b00101101; // Expected: {'P': 3195}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000111; B = 8'b00101101; | Outputs: P=%b | Expected: P=%d",
                 1387,
                 
                 P
                 , 
                 
                 3195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001110; B = 8'b01110101; // Expected: {'P': 24102}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001110; B = 8'b01110101; | Outputs: P=%b | Expected: P=%d",
                 1388,
                 
                 P
                 , 
                 
                 24102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000000; B = 8'b00010001; // Expected: {'P': 3264}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000000; B = 8'b00010001; | Outputs: P=%b | Expected: P=%d",
                 1389,
                 
                 P
                 , 
                 
                 3264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010111; B = 8'b00111011; // Expected: {'P': 1357}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010111; B = 8'b00111011; | Outputs: P=%b | Expected: P=%d",
                 1390,
                 
                 P
                 , 
                 
                 1357
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110001; B = 8'b00101111; // Expected: {'P': 8319}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110001; B = 8'b00101111; | Outputs: P=%b | Expected: P=%d",
                 1391,
                 
                 P
                 , 
                 
                 8319
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011100; B = 8'b00111100; // Expected: {'P': 13200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011100; B = 8'b00111100; | Outputs: P=%b | Expected: P=%d",
                 1392,
                 
                 P
                 , 
                 
                 13200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100111; B = 8'b10010100; // Expected: {'P': 15244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100111; B = 8'b10010100; | Outputs: P=%b | Expected: P=%d",
                 1393,
                 
                 P
                 , 
                 
                 15244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111101; B = 8'b01111010; // Expected: {'P': 23058}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111101; B = 8'b01111010; | Outputs: P=%b | Expected: P=%d",
                 1394,
                 
                 P
                 , 
                 
                 23058
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111001; B = 8'b00111100; // Expected: {'P': 7260}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111001; B = 8'b00111100; | Outputs: P=%b | Expected: P=%d",
                 1395,
                 
                 P
                 , 
                 
                 7260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010001; B = 8'b10001100; // Expected: {'P': 11340}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010001; B = 8'b10001100; | Outputs: P=%b | Expected: P=%d",
                 1396,
                 
                 P
                 , 
                 
                 11340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000100; B = 8'b10111000; // Expected: {'P': 736}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000100; B = 8'b10111000; | Outputs: P=%b | Expected: P=%d",
                 1397,
                 
                 P
                 , 
                 
                 736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011100; B = 8'b10011000; // Expected: {'P': 33440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011100; B = 8'b10011000; | Outputs: P=%b | Expected: P=%d",
                 1398,
                 
                 P
                 , 
                 
                 33440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101000; B = 8'b11000111; // Expected: {'P': 20696}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101000; B = 8'b11000111; | Outputs: P=%b | Expected: P=%d",
                 1399,
                 
                 P
                 , 
                 
                 20696
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111011; B = 8'b00001000; // Expected: {'P': 984}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111011; B = 8'b00001000; | Outputs: P=%b | Expected: P=%d",
                 1400,
                 
                 P
                 , 
                 
                 984
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010100; B = 8'b10101001; // Expected: {'P': 14196}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010100; B = 8'b10101001; | Outputs: P=%b | Expected: P=%d",
                 1401,
                 
                 P
                 , 
                 
                 14196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001011; B = 8'b10011001; // Expected: {'P': 11475}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001011; B = 8'b10011001; | Outputs: P=%b | Expected: P=%d",
                 1402,
                 
                 P
                 , 
                 
                 11475
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010110; B = 8'b10100000; // Expected: {'P': 3520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010110; B = 8'b10100000; | Outputs: P=%b | Expected: P=%d",
                 1403,
                 
                 P
                 , 
                 
                 3520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100111; B = 8'b10111111; // Expected: {'P': 7449}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100111; B = 8'b10111111; | Outputs: P=%b | Expected: P=%d",
                 1404,
                 
                 P
                 , 
                 
                 7449
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111010; B = 8'b11100100; // Expected: {'P': 13224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111010; B = 8'b11100100; | Outputs: P=%b | Expected: P=%d",
                 1405,
                 
                 P
                 , 
                 
                 13224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101010; B = 8'b01100111; // Expected: {'P': 17510}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101010; B = 8'b01100111; | Outputs: P=%b | Expected: P=%d",
                 1406,
                 
                 P
                 , 
                 
                 17510
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110111; B = 8'b10001011; // Expected: {'P': 7645}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110111; B = 8'b10001011; | Outputs: P=%b | Expected: P=%d",
                 1407,
                 
                 P
                 , 
                 
                 7645
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100111; B = 8'b11010001; // Expected: {'P': 21527}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100111; B = 8'b11010001; | Outputs: P=%b | Expected: P=%d",
                 1408,
                 
                 P
                 , 
                 
                 21527
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011000; B = 8'b10110110; // Expected: {'P': 39312}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011000; B = 8'b10110110; | Outputs: P=%b | Expected: P=%d",
                 1409,
                 
                 P
                 , 
                 
                 39312
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011111; B = 8'b01010101; // Expected: {'P': 8075}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011111; B = 8'b01010101; | Outputs: P=%b | Expected: P=%d",
                 1410,
                 
                 P
                 , 
                 
                 8075
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101111; B = 8'b01110000; // Expected: {'P': 19600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101111; B = 8'b01110000; | Outputs: P=%b | Expected: P=%d",
                 1411,
                 
                 P
                 , 
                 
                 19600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000110; B = 8'b10001001; // Expected: {'P': 822}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000110; B = 8'b10001001; | Outputs: P=%b | Expected: P=%d",
                 1412,
                 
                 P
                 , 
                 
                 822
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011000; B = 8'b11110101; // Expected: {'P': 52920}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011000; B = 8'b11110101; | Outputs: P=%b | Expected: P=%d",
                 1413,
                 
                 P
                 , 
                 
                 52920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001100; B = 8'b00101110; // Expected: {'P': 552}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001100; B = 8'b00101110; | Outputs: P=%b | Expected: P=%d",
                 1414,
                 
                 P
                 , 
                 
                 552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011100; B = 8'b01100000; // Expected: {'P': 8832}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011100; B = 8'b01100000; | Outputs: P=%b | Expected: P=%d",
                 1415,
                 
                 P
                 , 
                 
                 8832
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111010; B = 8'b01011100; // Expected: {'P': 17112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111010; B = 8'b01011100; | Outputs: P=%b | Expected: P=%d",
                 1416,
                 
                 P
                 , 
                 
                 17112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100110; B = 8'b00110011; // Expected: {'P': 5202}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100110; B = 8'b00110011; | Outputs: P=%b | Expected: P=%d",
                 1417,
                 
                 P
                 , 
                 
                 5202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110111; B = 8'b10111001; // Expected: {'P': 33855}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110111; B = 8'b10111001; | Outputs: P=%b | Expected: P=%d",
                 1418,
                 
                 P
                 , 
                 
                 33855
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101101; B = 8'b11111011; // Expected: {'P': 27359}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101101; B = 8'b11111011; | Outputs: P=%b | Expected: P=%d",
                 1419,
                 
                 P
                 , 
                 
                 27359
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101100; B = 8'b10011110; // Expected: {'P': 17064}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101100; B = 8'b10011110; | Outputs: P=%b | Expected: P=%d",
                 1420,
                 
                 P
                 , 
                 
                 17064
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001111; B = 8'b11000000; // Expected: {'P': 39744}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001111; B = 8'b11000000; | Outputs: P=%b | Expected: P=%d",
                 1421,
                 
                 P
                 , 
                 
                 39744
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101101; B = 8'b11000100; // Expected: {'P': 21364}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101101; B = 8'b11000100; | Outputs: P=%b | Expected: P=%d",
                 1422,
                 
                 P
                 , 
                 
                 21364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111100; B = 8'b11100011; // Expected: {'P': 57204}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111100; B = 8'b11100011; | Outputs: P=%b | Expected: P=%d",
                 1423,
                 
                 P
                 , 
                 
                 57204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110110; B = 8'b10011010; // Expected: {'P': 28028}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110110; B = 8'b10011010; | Outputs: P=%b | Expected: P=%d",
                 1424,
                 
                 P
                 , 
                 
                 28028
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101000; B = 8'b10101011; // Expected: {'P': 6840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101000; B = 8'b10101011; | Outputs: P=%b | Expected: P=%d",
                 1425,
                 
                 P
                 , 
                 
                 6840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001010; B = 8'b00000010; // Expected: {'P': 404}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001010; B = 8'b00000010; | Outputs: P=%b | Expected: P=%d",
                 1426,
                 
                 P
                 , 
                 
                 404
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110111; B = 8'b11101111; // Expected: {'P': 28441}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110111; B = 8'b11101111; | Outputs: P=%b | Expected: P=%d",
                 1427,
                 
                 P
                 , 
                 
                 28441
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000101; B = 8'b01001001; // Expected: {'P': 5037}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000101; B = 8'b01001001; | Outputs: P=%b | Expected: P=%d",
                 1428,
                 
                 P
                 , 
                 
                 5037
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010010; B = 8'b00101100; // Expected: {'P': 6424}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010010; B = 8'b00101100; | Outputs: P=%b | Expected: P=%d",
                 1429,
                 
                 P
                 , 
                 
                 6424
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000001; B = 8'b10100011; // Expected: {'P': 163}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000001; B = 8'b10100011; | Outputs: P=%b | Expected: P=%d",
                 1430,
                 
                 P
                 , 
                 
                 163
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111110; B = 8'b01010101; // Expected: {'P': 21590}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111110; B = 8'b01010101; | Outputs: P=%b | Expected: P=%d",
                 1431,
                 
                 P
                 , 
                 
                 21590
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011001; B = 8'b10100101; // Expected: {'P': 14685}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011001; B = 8'b10100101; | Outputs: P=%b | Expected: P=%d",
                 1432,
                 
                 P
                 , 
                 
                 14685
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101001; B = 8'b01001011; // Expected: {'P': 12675}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101001; B = 8'b01001011; | Outputs: P=%b | Expected: P=%d",
                 1433,
                 
                 P
                 , 
                 
                 12675
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010010; B = 8'b00011111; // Expected: {'P': 558}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010010; B = 8'b00011111; | Outputs: P=%b | Expected: P=%d",
                 1434,
                 
                 P
                 , 
                 
                 558
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001111; B = 8'b00111011; // Expected: {'P': 885}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001111; B = 8'b00111011; | Outputs: P=%b | Expected: P=%d",
                 1435,
                 
                 P
                 , 
                 
                 885
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100111; B = 8'b00100010; // Expected: {'P': 3502}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100111; B = 8'b00100010; | Outputs: P=%b | Expected: P=%d",
                 1436,
                 
                 P
                 , 
                 
                 3502
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001011; B = 8'b11111011; // Expected: {'P': 18825}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001011; B = 8'b11111011; | Outputs: P=%b | Expected: P=%d",
                 1437,
                 
                 P
                 , 
                 
                 18825
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010110; B = 8'b11010011; // Expected: {'P': 45154}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010110; B = 8'b11010011; | Outputs: P=%b | Expected: P=%d",
                 1438,
                 
                 P
                 , 
                 
                 45154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011000; B = 8'b10001011; // Expected: {'P': 30024}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011000; B = 8'b10001011; | Outputs: P=%b | Expected: P=%d",
                 1439,
                 
                 P
                 , 
                 
                 30024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110000; B = 8'b00010001; // Expected: {'P': 2992}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110000; B = 8'b00010001; | Outputs: P=%b | Expected: P=%d",
                 1440,
                 
                 P
                 , 
                 
                 2992
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100111; B = 8'b10000010; // Expected: {'P': 5070}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100111; B = 8'b10000010; | Outputs: P=%b | Expected: P=%d",
                 1441,
                 
                 P
                 , 
                 
                 5070
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111011; B = 8'b11001010; // Expected: {'P': 11918}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111011; B = 8'b11001010; | Outputs: P=%b | Expected: P=%d",
                 1442,
                 
                 P
                 , 
                 
                 11918
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011010; B = 8'b00000101; // Expected: {'P': 770}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011010; B = 8'b00000101; | Outputs: P=%b | Expected: P=%d",
                 1443,
                 
                 P
                 , 
                 
                 770
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100000; B = 8'b00101011; // Expected: {'P': 1376}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100000; B = 8'b00101011; | Outputs: P=%b | Expected: P=%d",
                 1444,
                 
                 P
                 , 
                 
                 1376
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000111; B = 8'b11011001; // Expected: {'P': 15407}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000111; B = 8'b11011001; | Outputs: P=%b | Expected: P=%d",
                 1445,
                 
                 P
                 , 
                 
                 15407
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011011; B = 8'b00111110; // Expected: {'P': 5642}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011011; B = 8'b00111110; | Outputs: P=%b | Expected: P=%d",
                 1446,
                 
                 P
                 , 
                 
                 5642
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100010; B = 8'b10011000; // Expected: {'P': 14896}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100010; B = 8'b10011000; | Outputs: P=%b | Expected: P=%d",
                 1447,
                 
                 P
                 , 
                 
                 14896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101110; B = 8'b10110101; // Expected: {'P': 8326}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101110; B = 8'b10110101; | Outputs: P=%b | Expected: P=%d",
                 1448,
                 
                 P
                 , 
                 
                 8326
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111000; B = 8'b10100100; // Expected: {'P': 19680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111000; B = 8'b10100100; | Outputs: P=%b | Expected: P=%d",
                 1449,
                 
                 P
                 , 
                 
                 19680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110111; B = 8'b11110010; // Expected: {'P': 59774}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110111; B = 8'b11110010; | Outputs: P=%b | Expected: P=%d",
                 1450,
                 
                 P
                 , 
                 
                 59774
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110111; B = 8'b00100010; // Expected: {'P': 4046}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110111; B = 8'b00100010; | Outputs: P=%b | Expected: P=%d",
                 1451,
                 
                 P
                 , 
                 
                 4046
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100100; B = 8'b01000011; // Expected: {'P': 2412}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100100; B = 8'b01000011; | Outputs: P=%b | Expected: P=%d",
                 1452,
                 
                 P
                 , 
                 
                 2412
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000111; B = 8'b01101100; // Expected: {'P': 756}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000111; B = 8'b01101100; | Outputs: P=%b | Expected: P=%d",
                 1453,
                 
                 P
                 , 
                 
                 756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100001; B = 8'b10000000; // Expected: {'P': 12416}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100001; B = 8'b10000000; | Outputs: P=%b | Expected: P=%d",
                 1454,
                 
                 P
                 , 
                 
                 12416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101011; B = 8'b11101010; // Expected: {'P': 54990}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101011; B = 8'b11101010; | Outputs: P=%b | Expected: P=%d",
                 1455,
                 
                 P
                 , 
                 
                 54990
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000010; B = 8'b11011100; // Expected: {'P': 28600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000010; B = 8'b11011100; | Outputs: P=%b | Expected: P=%d",
                 1456,
                 
                 P
                 , 
                 
                 28600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111111; B = 8'b11010000; // Expected: {'P': 13104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111111; B = 8'b11010000; | Outputs: P=%b | Expected: P=%d",
                 1457,
                 
                 P
                 , 
                 
                 13104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100011; B = 8'b01011010; // Expected: {'P': 8910}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100011; B = 8'b01011010; | Outputs: P=%b | Expected: P=%d",
                 1458,
                 
                 P
                 , 
                 
                 8910
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000100; B = 8'b10100000; // Expected: {'P': 31360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000100; B = 8'b10100000; | Outputs: P=%b | Expected: P=%d",
                 1459,
                 
                 P
                 , 
                 
                 31360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010110; B = 8'b10111101; // Expected: {'P': 16254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010110; B = 8'b10111101; | Outputs: P=%b | Expected: P=%d",
                 1460,
                 
                 P
                 , 
                 
                 16254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000111; B = 8'b10100010; // Expected: {'P': 32238}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000111; B = 8'b10100010; | Outputs: P=%b | Expected: P=%d",
                 1461,
                 
                 P
                 , 
                 
                 32238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111111; B = 8'b11011110; // Expected: {'P': 56610}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111111; B = 8'b11011110; | Outputs: P=%b | Expected: P=%d",
                 1462,
                 
                 P
                 , 
                 
                 56610
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000001; B = 8'b01001001; // Expected: {'P': 9417}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000001; B = 8'b01001001; | Outputs: P=%b | Expected: P=%d",
                 1463,
                 
                 P
                 , 
                 
                 9417
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000101; B = 8'b11111010; // Expected: {'P': 49250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000101; B = 8'b11111010; | Outputs: P=%b | Expected: P=%d",
                 1464,
                 
                 P
                 , 
                 
                 49250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010101; B = 8'b10101111; // Expected: {'P': 3675}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010101; B = 8'b10101111; | Outputs: P=%b | Expected: P=%d",
                 1465,
                 
                 P
                 , 
                 
                 3675
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001100; B = 8'b00011000; // Expected: {'P': 4896}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001100; B = 8'b00011000; | Outputs: P=%b | Expected: P=%d",
                 1466,
                 
                 P
                 , 
                 
                 4896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001001; B = 8'b01001001; // Expected: {'P': 10001}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001001; B = 8'b01001001; | Outputs: P=%b | Expected: P=%d",
                 1467,
                 
                 P
                 , 
                 
                 10001
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000100; B = 8'b00001101; // Expected: {'P': 1716}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000100; B = 8'b00001101; | Outputs: P=%b | Expected: P=%d",
                 1468,
                 
                 P
                 , 
                 
                 1716
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100001; B = 8'b10110011; // Expected: {'P': 28819}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100001; B = 8'b10110011; | Outputs: P=%b | Expected: P=%d",
                 1469,
                 
                 P
                 , 
                 
                 28819
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111011; B = 8'b00100001; // Expected: {'P': 4059}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111011; B = 8'b00100001; | Outputs: P=%b | Expected: P=%d",
                 1470,
                 
                 P
                 , 
                 
                 4059
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100001; B = 8'b10000101; // Expected: {'P': 29925}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100001; B = 8'b10000101; | Outputs: P=%b | Expected: P=%d",
                 1471,
                 
                 P
                 , 
                 
                 29925
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010001; B = 8'b10101000; // Expected: {'P': 2856}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010001; B = 8'b10101000; | Outputs: P=%b | Expected: P=%d",
                 1472,
                 
                 P
                 , 
                 
                 2856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011100; B = 8'b10100111; // Expected: {'P': 26052}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011100; B = 8'b10100111; | Outputs: P=%b | Expected: P=%d",
                 1473,
                 
                 P
                 , 
                 
                 26052
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001010; B = 8'b11011101; // Expected: {'P': 2210}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001010; B = 8'b11011101; | Outputs: P=%b | Expected: P=%d",
                 1474,
                 
                 P
                 , 
                 
                 2210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101101; B = 8'b10000010; // Expected: {'P': 22490}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101101; B = 8'b10000010; | Outputs: P=%b | Expected: P=%d",
                 1475,
                 
                 P
                 , 
                 
                 22490
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101101; B = 8'b11101010; // Expected: {'P': 55458}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101101; B = 8'b11101010; | Outputs: P=%b | Expected: P=%d",
                 1476,
                 
                 P
                 , 
                 
                 55458
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111001; B = 8'b01111111; // Expected: {'P': 23495}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111001; B = 8'b01111111; | Outputs: P=%b | Expected: P=%d",
                 1477,
                 
                 P
                 , 
                 
                 23495
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110101; B = 8'b00110111; // Expected: {'P': 6435}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110101; B = 8'b00110111; | Outputs: P=%b | Expected: P=%d",
                 1478,
                 
                 P
                 , 
                 
                 6435
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111101; B = 8'b00000111; // Expected: {'P': 1323}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111101; B = 8'b00000111; | Outputs: P=%b | Expected: P=%d",
                 1479,
                 
                 P
                 , 
                 
                 1323
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100001; B = 8'b11100101; // Expected: {'P': 36869}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100001; B = 8'b11100101; | Outputs: P=%b | Expected: P=%d",
                 1480,
                 
                 P
                 , 
                 
                 36869
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010011; B = 8'b11011111; // Expected: {'P': 32781}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010011; B = 8'b11011111; | Outputs: P=%b | Expected: P=%d",
                 1481,
                 
                 P
                 , 
                 
                 32781
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101100; B = 8'b01011010; // Expected: {'P': 21240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101100; B = 8'b01011010; | Outputs: P=%b | Expected: P=%d",
                 1482,
                 
                 P
                 , 
                 
                 21240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011110; B = 8'b10111110; // Expected: {'P': 5700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011110; B = 8'b10111110; | Outputs: P=%b | Expected: P=%d",
                 1483,
                 
                 P
                 , 
                 
                 5700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100100; B = 8'b11100000; // Expected: {'P': 51072}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100100; B = 8'b11100000; | Outputs: P=%b | Expected: P=%d",
                 1484,
                 
                 P
                 , 
                 
                 51072
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001100; B = 8'b11100011; // Expected: {'P': 31780}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001100; B = 8'b11100011; | Outputs: P=%b | Expected: P=%d",
                 1485,
                 
                 P
                 , 
                 
                 31780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100101; B = 8'b10010010; // Expected: {'P': 24090}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100101; B = 8'b10010010; | Outputs: P=%b | Expected: P=%d",
                 1486,
                 
                 P
                 , 
                 
                 24090
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011111; B = 8'b01001010; // Expected: {'P': 16502}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011111; B = 8'b01001010; | Outputs: P=%b | Expected: P=%d",
                 1487,
                 
                 P
                 , 
                 
                 16502
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101110; B = 8'b00110110; // Expected: {'P': 9396}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101110; B = 8'b00110110; | Outputs: P=%b | Expected: P=%d",
                 1488,
                 
                 P
                 , 
                 
                 9396
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011010; B = 8'b11000101; // Expected: {'P': 30338}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011010; B = 8'b11000101; | Outputs: P=%b | Expected: P=%d",
                 1489,
                 
                 P
                 , 
                 
                 30338
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111011; B = 8'b11010101; // Expected: {'P': 26199}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111011; B = 8'b11010101; | Outputs: P=%b | Expected: P=%d",
                 1490,
                 
                 P
                 , 
                 
                 26199
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101101; B = 8'b00101000; // Expected: {'P': 4360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101101; B = 8'b00101000; | Outputs: P=%b | Expected: P=%d",
                 1491,
                 
                 P
                 , 
                 
                 4360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100001; B = 8'b00011001; // Expected: {'P': 5625}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100001; B = 8'b00011001; | Outputs: P=%b | Expected: P=%d",
                 1492,
                 
                 P
                 , 
                 
                 5625
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000110; B = 8'b00110100; // Expected: {'P': 6968}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000110; B = 8'b00110100; | Outputs: P=%b | Expected: P=%d",
                 1493,
                 
                 P
                 , 
                 
                 6968
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011110; B = 8'b01000010; // Expected: {'P': 10428}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011110; B = 8'b01000010; | Outputs: P=%b | Expected: P=%d",
                 1494,
                 
                 P
                 , 
                 
                 10428
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000101; B = 8'b10111011; // Expected: {'P': 12903}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000101; B = 8'b10111011; | Outputs: P=%b | Expected: P=%d",
                 1495,
                 
                 P
                 , 
                 
                 12903
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001110; B = 8'b11011101; // Expected: {'P': 3094}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001110; B = 8'b11011101; | Outputs: P=%b | Expected: P=%d",
                 1496,
                 
                 P
                 , 
                 
                 3094
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011101; B = 8'b10101011; // Expected: {'P': 37791}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011101; B = 8'b10101011; | Outputs: P=%b | Expected: P=%d",
                 1497,
                 
                 P
                 , 
                 
                 37791
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110111; B = 8'b01000101; // Expected: {'P': 17043}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110111; B = 8'b01000101; | Outputs: P=%b | Expected: P=%d",
                 1498,
                 
                 P
                 , 
                 
                 17043
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101100; B = 8'b10100010; // Expected: {'P': 38232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101100; B = 8'b10100010; | Outputs: P=%b | Expected: P=%d",
                 1499,
                 
                 P
                 , 
                 
                 38232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010000; B = 8'b00010101; // Expected: {'P': 4368}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010000; B = 8'b00010101; | Outputs: P=%b | Expected: P=%d",
                 1500,
                 
                 P
                 , 
                 
                 4368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100000; B = 8'b11010011; // Expected: {'P': 20256}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100000; B = 8'b11010011; | Outputs: P=%b | Expected: P=%d",
                 1501,
                 
                 P
                 , 
                 
                 20256
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010010; B = 8'b11011011; // Expected: {'P': 31974}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010010; B = 8'b11011011; | Outputs: P=%b | Expected: P=%d",
                 1502,
                 
                 P
                 , 
                 
                 31974
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011110; B = 8'b01010010; // Expected: {'P': 18204}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011110; B = 8'b01010010; | Outputs: P=%b | Expected: P=%d",
                 1503,
                 
                 P
                 , 
                 
                 18204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111011; B = 8'b01110101; // Expected: {'P': 29367}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111011; B = 8'b01110101; | Outputs: P=%b | Expected: P=%d",
                 1504,
                 
                 P
                 , 
                 
                 29367
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110011; B = 8'b10100100; // Expected: {'P': 39852}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110011; B = 8'b10100100; | Outputs: P=%b | Expected: P=%d",
                 1505,
                 
                 P
                 , 
                 
                 39852
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100110; B = 8'b01010001; // Expected: {'P': 8262}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100110; B = 8'b01010001; | Outputs: P=%b | Expected: P=%d",
                 1506,
                 
                 P
                 , 
                 
                 8262
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010101; B = 8'b10100011; // Expected: {'P': 3423}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010101; B = 8'b10100011; | Outputs: P=%b | Expected: P=%d",
                 1507,
                 
                 P
                 , 
                 
                 3423
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001001; B = 8'b00101111; // Expected: {'P': 423}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001001; B = 8'b00101111; | Outputs: P=%b | Expected: P=%d",
                 1508,
                 
                 P
                 , 
                 
                 423
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001011; B = 8'b10011110; // Expected: {'P': 1738}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001011; B = 8'b10011110; | Outputs: P=%b | Expected: P=%d",
                 1509,
                 
                 P
                 , 
                 
                 1738
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100010; B = 8'b01011000; // Expected: {'P': 14256}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100010; B = 8'b01011000; | Outputs: P=%b | Expected: P=%d",
                 1510,
                 
                 P
                 , 
                 
                 14256
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000010; B = 8'b10011010; // Expected: {'P': 29876}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000010; B = 8'b10011010; | Outputs: P=%b | Expected: P=%d",
                 1511,
                 
                 P
                 , 
                 
                 29876
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011001; B = 8'b10000111; // Expected: {'P': 20655}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011001; B = 8'b10000111; | Outputs: P=%b | Expected: P=%d",
                 1512,
                 
                 P
                 , 
                 
                 20655
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010110; B = 8'b10001001; // Expected: {'P': 3014}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010110; B = 8'b10001001; | Outputs: P=%b | Expected: P=%d",
                 1513,
                 
                 P
                 , 
                 
                 3014
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001000; B = 8'b10111011; // Expected: {'P': 37400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001000; B = 8'b10111011; | Outputs: P=%b | Expected: P=%d",
                 1514,
                 
                 P
                 , 
                 
                 37400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111110; B = 8'b01001111; // Expected: {'P': 4898}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111110; B = 8'b01001111; | Outputs: P=%b | Expected: P=%d",
                 1515,
                 
                 P
                 , 
                 
                 4898
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011101; B = 8'b00011001; // Expected: {'P': 3925}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011101; B = 8'b00011001; | Outputs: P=%b | Expected: P=%d",
                 1516,
                 
                 P
                 , 
                 
                 3925
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110111; B = 8'b00111100; // Expected: {'P': 7140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110111; B = 8'b00111100; | Outputs: P=%b | Expected: P=%d",
                 1517,
                 
                 P
                 , 
                 
                 7140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101101; B = 8'b10100101; // Expected: {'P': 39105}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101101; B = 8'b10100101; | Outputs: P=%b | Expected: P=%d",
                 1518,
                 
                 P
                 , 
                 
                 39105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011101; B = 8'b01111101; // Expected: {'P': 27625}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011101; B = 8'b01111101; | Outputs: P=%b | Expected: P=%d",
                 1519,
                 
                 P
                 , 
                 
                 27625
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010100; B = 8'b10000110; // Expected: {'P': 2680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010100; B = 8'b10000110; | Outputs: P=%b | Expected: P=%d",
                 1520,
                 
                 P
                 , 
                 
                 2680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000011; B = 8'b01100011; // Expected: {'P': 297}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000011; B = 8'b01100011; | Outputs: P=%b | Expected: P=%d",
                 1521,
                 
                 P
                 , 
                 
                 297
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111100; B = 8'b00110110; // Expected: {'P': 3240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111100; B = 8'b00110110; | Outputs: P=%b | Expected: P=%d",
                 1522,
                 
                 P
                 , 
                 
                 3240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100001; B = 8'b00011000; // Expected: {'P': 2328}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100001; B = 8'b00011000; | Outputs: P=%b | Expected: P=%d",
                 1523,
                 
                 P
                 , 
                 
                 2328
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001010; B = 8'b10001000; // Expected: {'P': 18768}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001010; B = 8'b10001000; | Outputs: P=%b | Expected: P=%d",
                 1524,
                 
                 P
                 , 
                 
                 18768
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101010; B = 8'b10000011; // Expected: {'P': 5502}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101010; B = 8'b10000011; | Outputs: P=%b | Expected: P=%d",
                 1525,
                 
                 P
                 , 
                 
                 5502
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011111; B = 8'b10110000; // Expected: {'P': 5456}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011111; B = 8'b10110000; | Outputs: P=%b | Expected: P=%d",
                 1526,
                 
                 P
                 , 
                 
                 5456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000100; B = 8'b10100110; // Expected: {'P': 21912}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000100; B = 8'b10100110; | Outputs: P=%b | Expected: P=%d",
                 1527,
                 
                 P
                 , 
                 
                 21912
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110000; B = 8'b01001011; // Expected: {'P': 8400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110000; B = 8'b01001011; | Outputs: P=%b | Expected: P=%d",
                 1528,
                 
                 P
                 , 
                 
                 8400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000100; B = 8'b11011001; // Expected: {'P': 14756}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000100; B = 8'b11011001; | Outputs: P=%b | Expected: P=%d",
                 1529,
                 
                 P
                 , 
                 
                 14756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010001; B = 8'b00001000; // Expected: {'P': 1672}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010001; B = 8'b00001000; | Outputs: P=%b | Expected: P=%d",
                 1530,
                 
                 P
                 , 
                 
                 1672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110100; B = 8'b01011100; // Expected: {'P': 16560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110100; B = 8'b01011100; | Outputs: P=%b | Expected: P=%d",
                 1531,
                 
                 P
                 , 
                 
                 16560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110001; B = 8'b11110111; // Expected: {'P': 59527}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110001; B = 8'b11110111; | Outputs: P=%b | Expected: P=%d",
                 1532,
                 
                 P
                 , 
                 
                 59527
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111011; B = 8'b10011100; // Expected: {'P': 19188}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111011; B = 8'b10011100; | Outputs: P=%b | Expected: P=%d",
                 1533,
                 
                 P
                 , 
                 
                 19188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100111; B = 8'b10001011; // Expected: {'P': 14317}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100111; B = 8'b10001011; | Outputs: P=%b | Expected: P=%d",
                 1534,
                 
                 P
                 , 
                 
                 14317
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100110; B = 8'b01011101; // Expected: {'P': 3534}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100110; B = 8'b01011101; | Outputs: P=%b | Expected: P=%d",
                 1535,
                 
                 P
                 , 
                 
                 3534
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111000; B = 8'b11010000; // Expected: {'P': 51584}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111000; B = 8'b11010000; | Outputs: P=%b | Expected: P=%d",
                 1536,
                 
                 P
                 , 
                 
                 51584
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001001; B = 8'b10101110; // Expected: {'P': 12702}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001001; B = 8'b10101110; | Outputs: P=%b | Expected: P=%d",
                 1537,
                 
                 P
                 , 
                 
                 12702
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100011; B = 8'b10000001; // Expected: {'P': 12771}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100011; B = 8'b10000001; | Outputs: P=%b | Expected: P=%d",
                 1538,
                 
                 P
                 , 
                 
                 12771
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110110; B = 8'b01110101; // Expected: {'P': 21294}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110110; B = 8'b01110101; | Outputs: P=%b | Expected: P=%d",
                 1539,
                 
                 P
                 , 
                 
                 21294
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011101; B = 8'b10010111; // Expected: {'P': 33371}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011101; B = 8'b10010111; | Outputs: P=%b | Expected: P=%d",
                 1540,
                 
                 P
                 , 
                 
                 33371
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101000; B = 8'b01101010; // Expected: {'P': 24592}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101000; B = 8'b01101010; | Outputs: P=%b | Expected: P=%d",
                 1541,
                 
                 P
                 , 
                 
                 24592
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000010; B = 8'b11000000; // Expected: {'P': 24960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000010; B = 8'b11000000; | Outputs: P=%b | Expected: P=%d",
                 1542,
                 
                 P
                 , 
                 
                 24960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111100; B = 8'b01000110; // Expected: {'P': 17640}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111100; B = 8'b01000110; | Outputs: P=%b | Expected: P=%d",
                 1543,
                 
                 P
                 , 
                 
                 17640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001001; B = 8'b01100001; // Expected: {'P': 19497}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001001; B = 8'b01100001; | Outputs: P=%b | Expected: P=%d",
                 1544,
                 
                 P
                 , 
                 
                 19497
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011011; B = 8'b01101101; // Expected: {'P': 9919}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011011; B = 8'b01101101; | Outputs: P=%b | Expected: P=%d",
                 1545,
                 
                 P
                 , 
                 
                 9919
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111100; B = 8'b00111110; // Expected: {'P': 7688}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111100; B = 8'b00111110; | Outputs: P=%b | Expected: P=%d",
                 1546,
                 
                 P
                 , 
                 
                 7688
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010101; B = 8'b11010111; // Expected: {'P': 18275}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010101; B = 8'b11010111; | Outputs: P=%b | Expected: P=%d",
                 1547,
                 
                 P
                 , 
                 
                 18275
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101110; B = 8'b11111100; // Expected: {'P': 27720}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101110; B = 8'b11111100; | Outputs: P=%b | Expected: P=%d",
                 1548,
                 
                 P
                 , 
                 
                 27720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100100; B = 8'b11101101; // Expected: {'P': 8532}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100100; B = 8'b11101101; | Outputs: P=%b | Expected: P=%d",
                 1549,
                 
                 P
                 , 
                 
                 8532
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001000; B = 8'b10110011; // Expected: {'P': 35800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001000; B = 8'b10110011; | Outputs: P=%b | Expected: P=%d",
                 1550,
                 
                 P
                 , 
                 
                 35800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101100; B = 8'b00000111; // Expected: {'P': 1652}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101100; B = 8'b00000111; | Outputs: P=%b | Expected: P=%d",
                 1551,
                 
                 P
                 , 
                 
                 1652
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101010; B = 8'b10111001; // Expected: {'P': 7770}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101010; B = 8'b10111001; | Outputs: P=%b | Expected: P=%d",
                 1552,
                 
                 P
                 , 
                 
                 7770
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001000; B = 8'b10011100; // Expected: {'P': 11232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001000; B = 8'b10011100; | Outputs: P=%b | Expected: P=%d",
                 1553,
                 
                 P
                 , 
                 
                 11232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001010; B = 8'b11000000; // Expected: {'P': 14208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001010; B = 8'b11000000; | Outputs: P=%b | Expected: P=%d",
                 1554,
                 
                 P
                 , 
                 
                 14208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011001; B = 8'b11000000; // Expected: {'P': 17088}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011001; B = 8'b11000000; | Outputs: P=%b | Expected: P=%d",
                 1555,
                 
                 P
                 , 
                 
                 17088
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101111; B = 8'b10100101; // Expected: {'P': 39435}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101111; B = 8'b10100101; | Outputs: P=%b | Expected: P=%d",
                 1556,
                 
                 P
                 , 
                 
                 39435
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110101; B = 8'b11011100; // Expected: {'P': 25740}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110101; B = 8'b11011100; | Outputs: P=%b | Expected: P=%d",
                 1557,
                 
                 P
                 , 
                 
                 25740
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111101; B = 8'b01010111; // Expected: {'P': 5307}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111101; B = 8'b01010111; | Outputs: P=%b | Expected: P=%d",
                 1558,
                 
                 P
                 , 
                 
                 5307
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111101; B = 8'b11101101; // Expected: {'P': 14457}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111101; B = 8'b11101101; | Outputs: P=%b | Expected: P=%d",
                 1559,
                 
                 P
                 , 
                 
                 14457
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010001; B = 8'b01111100; // Expected: {'P': 10044}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010001; B = 8'b01111100; | Outputs: P=%b | Expected: P=%d",
                 1560,
                 
                 P
                 , 
                 
                 10044
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011110; B = 8'b10001000; // Expected: {'P': 4080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011110; B = 8'b10001000; | Outputs: P=%b | Expected: P=%d",
                 1561,
                 
                 P
                 , 
                 
                 4080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011000; B = 8'b00011001; // Expected: {'P': 2200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011000; B = 8'b00011001; | Outputs: P=%b | Expected: P=%d",
                 1562,
                 
                 P
                 , 
                 
                 2200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000101; B = 8'b11111001; // Expected: {'P': 1245}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000101; B = 8'b11111001; | Outputs: P=%b | Expected: P=%d",
                 1563,
                 
                 P
                 , 
                 
                 1245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001111; B = 8'b01110100; // Expected: {'P': 9164}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001111; B = 8'b01110100; | Outputs: P=%b | Expected: P=%d",
                 1564,
                 
                 P
                 , 
                 
                 9164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100101; B = 8'b10110100; // Expected: {'P': 6660}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100101; B = 8'b10110100; | Outputs: P=%b | Expected: P=%d",
                 1565,
                 
                 P
                 , 
                 
                 6660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011000; B = 8'b10111100; // Expected: {'P': 28576}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011000; B = 8'b10111100; | Outputs: P=%b | Expected: P=%d",
                 1566,
                 
                 P
                 , 
                 
                 28576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011101; B = 8'b11111101; // Expected: {'P': 23529}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011101; B = 8'b11111101; | Outputs: P=%b | Expected: P=%d",
                 1567,
                 
                 P
                 , 
                 
                 23529
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101001; B = 8'b10110110; // Expected: {'P': 42406}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101001; B = 8'b10110110; | Outputs: P=%b | Expected: P=%d",
                 1568,
                 
                 P
                 , 
                 
                 42406
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101101; B = 8'b11111100; // Expected: {'P': 43596}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101101; B = 8'b11111100; | Outputs: P=%b | Expected: P=%d",
                 1569,
                 
                 P
                 , 
                 
                 43596
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011011; B = 8'b10000000; // Expected: {'P': 19840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011011; B = 8'b10000000; | Outputs: P=%b | Expected: P=%d",
                 1570,
                 
                 P
                 , 
                 
                 19840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110111; B = 8'b01011111; // Expected: {'P': 23465}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110111; B = 8'b01011111; | Outputs: P=%b | Expected: P=%d",
                 1571,
                 
                 P
                 , 
                 
                 23465
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000000; B = 8'b00110011; // Expected: {'P': 9792}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000000; B = 8'b00110011; | Outputs: P=%b | Expected: P=%d",
                 1572,
                 
                 P
                 , 
                 
                 9792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011010; B = 8'b11000111; // Expected: {'P': 5174}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011010; B = 8'b11000111; | Outputs: P=%b | Expected: P=%d",
                 1573,
                 
                 P
                 , 
                 
                 5174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111001; B = 8'b01100111; // Expected: {'P': 19055}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111001; B = 8'b01100111; | Outputs: P=%b | Expected: P=%d",
                 1574,
                 
                 P
                 , 
                 
                 19055
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010000; B = 8'b00010000; // Expected: {'P': 256}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010000; B = 8'b00010000; | Outputs: P=%b | Expected: P=%d",
                 1575,
                 
                 P
                 , 
                 
                 256
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100001; B = 8'b11110101; // Expected: {'P': 55125}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100001; B = 8'b11110101; | Outputs: P=%b | Expected: P=%d",
                 1576,
                 
                 P
                 , 
                 
                 55125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011110; B = 8'b01100110; // Expected: {'P': 3060}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011110; B = 8'b01100110; | Outputs: P=%b | Expected: P=%d",
                 1577,
                 
                 P
                 , 
                 
                 3060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101000; B = 8'b00101010; // Expected: {'P': 4368}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101000; B = 8'b00101010; | Outputs: P=%b | Expected: P=%d",
                 1578,
                 
                 P
                 , 
                 
                 4368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101001; B = 8'b11011100; // Expected: {'P': 51260}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101001; B = 8'b11011100; | Outputs: P=%b | Expected: P=%d",
                 1579,
                 
                 P
                 , 
                 
                 51260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010000; B = 8'b00110000; // Expected: {'P': 9984}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010000; B = 8'b00110000; | Outputs: P=%b | Expected: P=%d",
                 1580,
                 
                 P
                 , 
                 
                 9984
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011011; B = 8'b01100011; // Expected: {'P': 2673}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011011; B = 8'b01100011; | Outputs: P=%b | Expected: P=%d",
                 1581,
                 
                 P
                 , 
                 
                 2673
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101100; B = 8'b10000100; // Expected: {'P': 14256}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101100; B = 8'b10000100; | Outputs: P=%b | Expected: P=%d",
                 1582,
                 
                 P
                 , 
                 
                 14256
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110011; B = 8'b00101111; // Expected: {'P': 5405}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110011; B = 8'b00101111; | Outputs: P=%b | Expected: P=%d",
                 1583,
                 
                 P
                 , 
                 
                 5405
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110010; B = 8'b00010111; // Expected: {'P': 4094}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110010; B = 8'b00010111; | Outputs: P=%b | Expected: P=%d",
                 1584,
                 
                 P
                 , 
                 
                 4094
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010110; B = 8'b10011110; // Expected: {'P': 13588}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010110; B = 8'b10011110; | Outputs: P=%b | Expected: P=%d",
                 1585,
                 
                 P
                 , 
                 
                 13588
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100001; B = 8'b00110000; // Expected: {'P': 10800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100001; B = 8'b00110000; | Outputs: P=%b | Expected: P=%d",
                 1586,
                 
                 P
                 , 
                 
                 10800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100100; B = 8'b11110001; // Expected: {'P': 39524}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100100; B = 8'b11110001; | Outputs: P=%b | Expected: P=%d",
                 1587,
                 
                 P
                 , 
                 
                 39524
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111111; B = 8'b10100101; // Expected: {'P': 10395}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111111; B = 8'b10100101; | Outputs: P=%b | Expected: P=%d",
                 1588,
                 
                 P
                 , 
                 
                 10395
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101000; B = 8'b00010100; // Expected: {'P': 4640}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101000; B = 8'b00010100; | Outputs: P=%b | Expected: P=%d",
                 1589,
                 
                 P
                 , 
                 
                 4640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111011; B = 8'b10010111; // Expected: {'P': 8909}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111011; B = 8'b10010111; | Outputs: P=%b | Expected: P=%d",
                 1590,
                 
                 P
                 , 
                 
                 8909
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110110; B = 8'b00001011; // Expected: {'P': 2706}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110110; B = 8'b00001011; | Outputs: P=%b | Expected: P=%d",
                 1591,
                 
                 P
                 , 
                 
                 2706
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011100; B = 8'b01111000; // Expected: {'P': 26400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011100; B = 8'b01111000; | Outputs: P=%b | Expected: P=%d",
                 1592,
                 
                 P
                 , 
                 
                 26400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111101; B = 8'b01010001; // Expected: {'P': 15309}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111101; B = 8'b01010001; | Outputs: P=%b | Expected: P=%d",
                 1593,
                 
                 P
                 , 
                 
                 15309
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000101; B = 8'b11001100; // Expected: {'P': 14076}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000101; B = 8'b11001100; | Outputs: P=%b | Expected: P=%d",
                 1594,
                 
                 P
                 , 
                 
                 14076
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100001; B = 8'b00101101; // Expected: {'P': 7245}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100001; B = 8'b00101101; | Outputs: P=%b | Expected: P=%d",
                 1595,
                 
                 P
                 , 
                 
                 7245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000011; B = 8'b10011110; // Expected: {'P': 20698}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000011; B = 8'b10011110; | Outputs: P=%b | Expected: P=%d",
                 1596,
                 
                 P
                 , 
                 
                 20698
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110101; B = 8'b10101010; // Expected: {'P': 9010}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110101; B = 8'b10101010; | Outputs: P=%b | Expected: P=%d",
                 1597,
                 
                 P
                 , 
                 
                 9010
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001011; B = 8'b10110101; // Expected: {'P': 13575}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001011; B = 8'b10110101; | Outputs: P=%b | Expected: P=%d",
                 1598,
                 
                 P
                 , 
                 
                 13575
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010100; B = 8'b01000111; // Expected: {'P': 10508}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010100; B = 8'b01000111; | Outputs: P=%b | Expected: P=%d",
                 1599,
                 
                 P
                 , 
                 
                 10508
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100100; B = 8'b10111101; // Expected: {'P': 18900}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100100; B = 8'b10111101; | Outputs: P=%b | Expected: P=%d",
                 1600,
                 
                 P
                 , 
                 
                 18900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000001; B = 8'b00000010; // Expected: {'P': 386}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000001; B = 8'b00000010; | Outputs: P=%b | Expected: P=%d",
                 1601,
                 
                 P
                 , 
                 
                 386
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100001; B = 8'b00000101; // Expected: {'P': 485}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100001; B = 8'b00000101; | Outputs: P=%b | Expected: P=%d",
                 1602,
                 
                 P
                 , 
                 
                 485
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010100; B = 8'b00000101; // Expected: {'P': 740}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010100; B = 8'b00000101; | Outputs: P=%b | Expected: P=%d",
                 1603,
                 
                 P
                 , 
                 
                 740
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101010; B = 8'b11001000; // Expected: {'P': 8400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101010; B = 8'b11001000; | Outputs: P=%b | Expected: P=%d",
                 1604,
                 
                 P
                 , 
                 
                 8400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001001; B = 8'b01001100; // Expected: {'P': 15276}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001001; B = 8'b01001100; | Outputs: P=%b | Expected: P=%d",
                 1605,
                 
                 P
                 , 
                 
                 15276
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010010; B = 8'b01001011; // Expected: {'P': 6150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010010; B = 8'b01001011; | Outputs: P=%b | Expected: P=%d",
                 1606,
                 
                 P
                 , 
                 
                 6150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111011; B = 8'b00110100; // Expected: {'P': 3068}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111011; B = 8'b00110100; | Outputs: P=%b | Expected: P=%d",
                 1607,
                 
                 P
                 , 
                 
                 3068
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110011; B = 8'b11101000; // Expected: {'P': 26680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110011; B = 8'b11101000; | Outputs: P=%b | Expected: P=%d",
                 1608,
                 
                 P
                 , 
                 
                 26680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000010; B = 8'b11100000; // Expected: {'P': 14784}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000010; B = 8'b11100000; | Outputs: P=%b | Expected: P=%d",
                 1609,
                 
                 P
                 , 
                 
                 14784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111010; B = 8'b11010100; // Expected: {'P': 53000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111010; B = 8'b11010100; | Outputs: P=%b | Expected: P=%d",
                 1610,
                 
                 P
                 , 
                 
                 53000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010010; B = 8'b01010101; // Expected: {'P': 6970}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010010; B = 8'b01010101; | Outputs: P=%b | Expected: P=%d",
                 1611,
                 
                 P
                 , 
                 
                 6970
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001110; B = 8'b00111100; // Expected: {'P': 8520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001110; B = 8'b00111100; | Outputs: P=%b | Expected: P=%d",
                 1612,
                 
                 P
                 , 
                 
                 8520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110101; B = 8'b01011110; // Expected: {'P': 10998}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110101; B = 8'b01011110; | Outputs: P=%b | Expected: P=%d",
                 1613,
                 
                 P
                 , 
                 
                 10998
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011101; B = 8'b10010100; // Expected: {'P': 13764}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011101; B = 8'b10010100; | Outputs: P=%b | Expected: P=%d",
                 1614,
                 
                 P
                 , 
                 
                 13764
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001011; B = 8'b00011101; // Expected: {'P': 2175}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001011; B = 8'b00011101; | Outputs: P=%b | Expected: P=%d",
                 1615,
                 
                 P
                 , 
                 
                 2175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001100; B = 8'b01001011; // Expected: {'P': 10500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001100; B = 8'b01001011; | Outputs: P=%b | Expected: P=%d",
                 1616,
                 
                 P
                 , 
                 
                 10500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110000; B = 8'b10011100; // Expected: {'P': 27456}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110000; B = 8'b10011100; | Outputs: P=%b | Expected: P=%d",
                 1617,
                 
                 P
                 , 
                 
                 27456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101110; B = 8'b11011111; // Expected: {'P': 53074}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101110; B = 8'b11011111; | Outputs: P=%b | Expected: P=%d",
                 1618,
                 
                 P
                 , 
                 
                 53074
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001010; B = 8'b00000110; // Expected: {'P': 1212}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001010; B = 8'b00000110; | Outputs: P=%b | Expected: P=%d",
                 1619,
                 
                 P
                 , 
                 
                 1212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010110; B = 8'b10110001; // Expected: {'P': 15222}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010110; B = 8'b10110001; | Outputs: P=%b | Expected: P=%d",
                 1620,
                 
                 P
                 , 
                 
                 15222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010000; B = 8'b10011111; // Expected: {'P': 12720}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010000; B = 8'b10011111; | Outputs: P=%b | Expected: P=%d",
                 1621,
                 
                 P
                 , 
                 
                 12720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101001; B = 8'b00001101; // Expected: {'P': 2197}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101001; B = 8'b00001101; | Outputs: P=%b | Expected: P=%d",
                 1622,
                 
                 P
                 , 
                 
                 2197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100100; B = 8'b10110101; // Expected: {'P': 6516}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100100; B = 8'b10110101; | Outputs: P=%b | Expected: P=%d",
                 1623,
                 
                 P
                 , 
                 
                 6516
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010101; B = 8'b10001100; // Expected: {'P': 2940}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010101; B = 8'b10001100; | Outputs: P=%b | Expected: P=%d",
                 1624,
                 
                 P
                 , 
                 
                 2940
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101101; B = 8'b11010100; // Expected: {'P': 23108}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101101; B = 8'b11010100; | Outputs: P=%b | Expected: P=%d",
                 1625,
                 
                 P
                 , 
                 
                 23108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110001; B = 8'b11011010; // Expected: {'P': 52538}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110001; B = 8'b11011010; | Outputs: P=%b | Expected: P=%d",
                 1626,
                 
                 P
                 , 
                 
                 52538
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100000; B = 8'b11110110; // Expected: {'P': 7872}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100000; B = 8'b11110110; | Outputs: P=%b | Expected: P=%d",
                 1627,
                 
                 P
                 , 
                 
                 7872
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000000; B = 8'b01011011; // Expected: {'P': 5824}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000000; B = 8'b01011011; | Outputs: P=%b | Expected: P=%d",
                 1628,
                 
                 P
                 , 
                 
                 5824
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001000; B = 8'b00010111; // Expected: {'P': 3128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001000; B = 8'b00010111; | Outputs: P=%b | Expected: P=%d",
                 1629,
                 
                 P
                 , 
                 
                 3128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100110; B = 8'b10101101; // Expected: {'P': 17646}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100110; B = 8'b10101101; | Outputs: P=%b | Expected: P=%d",
                 1630,
                 
                 P
                 , 
                 
                 17646
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110000; B = 8'b10111100; // Expected: {'P': 9024}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110000; B = 8'b10111100; | Outputs: P=%b | Expected: P=%d",
                 1631,
                 
                 P
                 , 
                 
                 9024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100011; B = 8'b11100111; // Expected: {'P': 52437}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100011; B = 8'b11100111; | Outputs: P=%b | Expected: P=%d",
                 1632,
                 
                 P
                 , 
                 
                 52437
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101110; B = 8'b11011101; // Expected: {'P': 10166}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101110; B = 8'b11011101; | Outputs: P=%b | Expected: P=%d",
                 1633,
                 
                 P
                 , 
                 
                 10166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001010; B = 8'b10110100; // Expected: {'P': 13320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001010; B = 8'b10110100; | Outputs: P=%b | Expected: P=%d",
                 1634,
                 
                 P
                 , 
                 
                 13320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011001; B = 8'b00010001; // Expected: {'P': 2601}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011001; B = 8'b00010001; | Outputs: P=%b | Expected: P=%d",
                 1635,
                 
                 P
                 , 
                 
                 2601
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011011; B = 8'b11111101; // Expected: {'P': 39215}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011011; B = 8'b11111101; | Outputs: P=%b | Expected: P=%d",
                 1636,
                 
                 P
                 , 
                 
                 39215
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000110; B = 8'b00111001; // Expected: {'P': 7638}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000110; B = 8'b00111001; | Outputs: P=%b | Expected: P=%d",
                 1637,
                 
                 P
                 , 
                 
                 7638
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110111; B = 8'b11110110; // Expected: {'P': 13530}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110111; B = 8'b11110110; | Outputs: P=%b | Expected: P=%d",
                 1638,
                 
                 P
                 , 
                 
                 13530
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100110; B = 8'b01111100; // Expected: {'P': 20584}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100110; B = 8'b01111100; | Outputs: P=%b | Expected: P=%d",
                 1639,
                 
                 P
                 , 
                 
                 20584
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110001; B = 8'b10100001; // Expected: {'P': 7889}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110001; B = 8'b10100001; | Outputs: P=%b | Expected: P=%d",
                 1640,
                 
                 P
                 , 
                 
                 7889
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110001; B = 8'b01110001; // Expected: {'P': 27233}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110001; B = 8'b01110001; | Outputs: P=%b | Expected: P=%d",
                 1641,
                 
                 P
                 , 
                 
                 27233
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011101; B = 8'b00001110; // Expected: {'P': 2198}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011101; B = 8'b00001110; | Outputs: P=%b | Expected: P=%d",
                 1642,
                 
                 P
                 , 
                 
                 2198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000011; B = 8'b11011001; // Expected: {'P': 14539}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000011; B = 8'b11011001; | Outputs: P=%b | Expected: P=%d",
                 1643,
                 
                 P
                 , 
                 
                 14539
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001100; B = 8'b10000000; // Expected: {'P': 26112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001100; B = 8'b10000000; | Outputs: P=%b | Expected: P=%d",
                 1644,
                 
                 P
                 , 
                 
                 26112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111100; B = 8'b01000000; // Expected: {'P': 3840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111100; B = 8'b01000000; | Outputs: P=%b | Expected: P=%d",
                 1645,
                 
                 P
                 , 
                 
                 3840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010101; B = 8'b11011001; // Expected: {'P': 4557}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010101; B = 8'b11011001; | Outputs: P=%b | Expected: P=%d",
                 1646,
                 
                 P
                 , 
                 
                 4557
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100110; B = 8'b10011100; // Expected: {'P': 25896}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100110; B = 8'b10011100; | Outputs: P=%b | Expected: P=%d",
                 1647,
                 
                 P
                 , 
                 
                 25896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111111; B = 8'b00000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111111; B = 8'b00000000; | Outputs: P=%b | Expected: P=%d",
                 1648,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001100; B = 8'b10110111; // Expected: {'P': 25620}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001100; B = 8'b10110111; | Outputs: P=%b | Expected: P=%d",
                 1649,
                 
                 P
                 , 
                 
                 25620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101010; B = 8'b01001011; // Expected: {'P': 7950}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101010; B = 8'b01001011; | Outputs: P=%b | Expected: P=%d",
                 1650,
                 
                 P
                 , 
                 
                 7950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001011; B = 8'b10001101; // Expected: {'P': 19599}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001011; B = 8'b10001101; | Outputs: P=%b | Expected: P=%d",
                 1651,
                 
                 P
                 , 
                 
                 19599
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111101; B = 8'b10000110; // Expected: {'P': 33902}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111101; B = 8'b10000110; | Outputs: P=%b | Expected: P=%d",
                 1652,
                 
                 P
                 , 
                 
                 33902
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010011; B = 8'b10111011; // Expected: {'P': 39457}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010011; B = 8'b10111011; | Outputs: P=%b | Expected: P=%d",
                 1653,
                 
                 P
                 , 
                 
                 39457
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110100; B = 8'b11100111; // Expected: {'P': 12012}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110100; B = 8'b11100111; | Outputs: P=%b | Expected: P=%d",
                 1654,
                 
                 P
                 , 
                 
                 12012
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101010; B = 8'b10001011; // Expected: {'P': 14734}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101010; B = 8'b10001011; | Outputs: P=%b | Expected: P=%d",
                 1655,
                 
                 P
                 , 
                 
                 14734
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001100; B = 8'b11010111; // Expected: {'P': 16340}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001100; B = 8'b11010111; | Outputs: P=%b | Expected: P=%d",
                 1656,
                 
                 P
                 , 
                 
                 16340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101011; B = 8'b10011011; // Expected: {'P': 6665}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101011; B = 8'b10011011; | Outputs: P=%b | Expected: P=%d",
                 1657,
                 
                 P
                 , 
                 
                 6665
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000111; B = 8'b00001011; // Expected: {'P': 1485}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000111; B = 8'b00001011; | Outputs: P=%b | Expected: P=%d",
                 1658,
                 
                 P
                 , 
                 
                 1485
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101010; B = 8'b00101011; // Expected: {'P': 7310}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101010; B = 8'b00101011; | Outputs: P=%b | Expected: P=%d",
                 1659,
                 
                 P
                 , 
                 
                 7310
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010110; B = 8'b01100101; // Expected: {'P': 21614}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010110; B = 8'b01100101; | Outputs: P=%b | Expected: P=%d",
                 1660,
                 
                 P
                 , 
                 
                 21614
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100101; B = 8'b11101111; // Expected: {'P': 24139}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100101; B = 8'b11101111; | Outputs: P=%b | Expected: P=%d",
                 1661,
                 
                 P
                 , 
                 
                 24139
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010011; B = 8'b10101000; // Expected: {'P': 3192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010011; B = 8'b10101000; | Outputs: P=%b | Expected: P=%d",
                 1662,
                 
                 P
                 , 
                 
                 3192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110010; B = 8'b10000111; // Expected: {'P': 32670}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110010; B = 8'b10000111; | Outputs: P=%b | Expected: P=%d",
                 1663,
                 
                 P
                 , 
                 
                 32670
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010001; B = 8'b01011001; // Expected: {'P': 12905}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010001; B = 8'b01011001; | Outputs: P=%b | Expected: P=%d",
                 1664,
                 
                 P
                 , 
                 
                 12905
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111010; B = 8'b11101101; // Expected: {'P': 44082}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111010; B = 8'b11101101; | Outputs: P=%b | Expected: P=%d",
                 1665,
                 
                 P
                 , 
                 
                 44082
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011101; B = 8'b11110111; // Expected: {'P': 38779}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011101; B = 8'b11110111; | Outputs: P=%b | Expected: P=%d",
                 1666,
                 
                 P
                 , 
                 
                 38779
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101001; B = 8'b01001110; // Expected: {'P': 8190}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101001; B = 8'b01001110; | Outputs: P=%b | Expected: P=%d",
                 1667,
                 
                 P
                 , 
                 
                 8190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101110; B = 8'b10110101; // Expected: {'P': 43078}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101110; B = 8'b10110101; | Outputs: P=%b | Expected: P=%d",
                 1668,
                 
                 P
                 , 
                 
                 43078
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011110; B = 8'b01000010; // Expected: {'P': 14652}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011110; B = 8'b01000010; | Outputs: P=%b | Expected: P=%d",
                 1669,
                 
                 P
                 , 
                 
                 14652
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010101; B = 8'b10100101; // Expected: {'P': 35145}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010101; B = 8'b10100101; | Outputs: P=%b | Expected: P=%d",
                 1670,
                 
                 P
                 , 
                 
                 35145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111101; B = 8'b10011100; // Expected: {'P': 9516}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111101; B = 8'b10011100; | Outputs: P=%b | Expected: P=%d",
                 1671,
                 
                 P
                 , 
                 
                 9516
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000001; B = 8'b11100101; // Expected: {'P': 29541}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000001; B = 8'b11100101; | Outputs: P=%b | Expected: P=%d",
                 1672,
                 
                 P
                 , 
                 
                 29541
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111101; B = 8'b10110110; // Expected: {'P': 46046}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111101; B = 8'b10110110; | Outputs: P=%b | Expected: P=%d",
                 1673,
                 
                 P
                 , 
                 
                 46046
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001000; B = 8'b11011101; // Expected: {'P': 1768}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001000; B = 8'b11011101; | Outputs: P=%b | Expected: P=%d",
                 1674,
                 
                 P
                 , 
                 
                 1768
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100001; B = 8'b10000110; // Expected: {'P': 4422}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100001; B = 8'b10000110; | Outputs: P=%b | Expected: P=%d",
                 1675,
                 
                 P
                 , 
                 
                 4422
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111111; B = 8'b00011001; // Expected: {'P': 1575}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111111; B = 8'b00011001; | Outputs: P=%b | Expected: P=%d",
                 1676,
                 
                 P
                 , 
                 
                 1575
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110010; B = 8'b01000101; // Expected: {'P': 16698}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110010; B = 8'b01000101; | Outputs: P=%b | Expected: P=%d",
                 1677,
                 
                 P
                 , 
                 
                 16698
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101000; B = 8'b01010101; // Expected: {'P': 8840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101000; B = 8'b01010101; | Outputs: P=%b | Expected: P=%d",
                 1678,
                 
                 P
                 , 
                 
                 8840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011000; B = 8'b00100010; // Expected: {'P': 5168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011000; B = 8'b00100010; | Outputs: P=%b | Expected: P=%d",
                 1679,
                 
                 P
                 , 
                 
                 5168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101111; B = 8'b10110100; // Expected: {'P': 19980}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101111; B = 8'b10110100; | Outputs: P=%b | Expected: P=%d",
                 1680,
                 
                 P
                 , 
                 
                 19980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111011; B = 8'b11001111; // Expected: {'P': 25461}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111011; B = 8'b11001111; | Outputs: P=%b | Expected: P=%d",
                 1681,
                 
                 P
                 , 
                 
                 25461
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100100; B = 8'b00110011; // Expected: {'P': 1836}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100100; B = 8'b00110011; | Outputs: P=%b | Expected: P=%d",
                 1682,
                 
                 P
                 , 
                 
                 1836
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101001; B = 8'b00100000; // Expected: {'P': 7456}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101001; B = 8'b00100000; | Outputs: P=%b | Expected: P=%d",
                 1683,
                 
                 P
                 , 
                 
                 7456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101000; B = 8'b11101001; // Expected: {'P': 9320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101000; B = 8'b11101001; | Outputs: P=%b | Expected: P=%d",
                 1684,
                 
                 P
                 , 
                 
                 9320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010010; B = 8'b00110010; // Expected: {'P': 7300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010010; B = 8'b00110010; | Outputs: P=%b | Expected: P=%d",
                 1685,
                 
                 P
                 , 
                 
                 7300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011001; B = 8'b10111110; // Expected: {'P': 4750}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011001; B = 8'b10111110; | Outputs: P=%b | Expected: P=%d",
                 1686,
                 
                 P
                 , 
                 
                 4750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110000; B = 8'b11101010; // Expected: {'P': 56160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110000; B = 8'b11101010; | Outputs: P=%b | Expected: P=%d",
                 1687,
                 
                 P
                 , 
                 
                 56160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010110; B = 8'b01010011; // Expected: {'P': 12450}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010110; B = 8'b01010011; | Outputs: P=%b | Expected: P=%d",
                 1688,
                 
                 P
                 , 
                 
                 12450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001001; B = 8'b01111110; // Expected: {'P': 1134}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001001; B = 8'b01111110; | Outputs: P=%b | Expected: P=%d",
                 1689,
                 
                 P
                 , 
                 
                 1134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010011; B = 8'b11011111; // Expected: {'P': 47053}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010011; B = 8'b11011111; | Outputs: P=%b | Expected: P=%d",
                 1690,
                 
                 P
                 , 
                 
                 47053
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010100; B = 8'b01111110; // Expected: {'P': 18648}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010100; B = 8'b01111110; | Outputs: P=%b | Expected: P=%d",
                 1691,
                 
                 P
                 , 
                 
                 18648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101010; B = 8'b01101011; // Expected: {'P': 25038}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101010; B = 8'b01101011; | Outputs: P=%b | Expected: P=%d",
                 1692,
                 
                 P
                 , 
                 
                 25038
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000101; B = 8'b11111010; // Expected: {'P': 1250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000101; B = 8'b11111010; | Outputs: P=%b | Expected: P=%d",
                 1693,
                 
                 P
                 , 
                 
                 1250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110111; B = 8'b10000000; // Expected: {'P': 7040}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110111; B = 8'b10000000; | Outputs: P=%b | Expected: P=%d",
                 1694,
                 
                 P
                 , 
                 
                 7040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101111; B = 8'b01001100; // Expected: {'P': 3572}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101111; B = 8'b01001100; | Outputs: P=%b | Expected: P=%d",
                 1695,
                 
                 P
                 , 
                 
                 3572
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101111; B = 8'b01110010; // Expected: {'P': 19950}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101111; B = 8'b01110010; | Outputs: P=%b | Expected: P=%d",
                 1696,
                 
                 P
                 , 
                 
                 19950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011110; B = 8'b00010101; // Expected: {'P': 1974}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011110; B = 8'b00010101; | Outputs: P=%b | Expected: P=%d",
                 1697,
                 
                 P
                 , 
                 
                 1974
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011011; B = 8'b01111110; // Expected: {'P': 27594}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011011; B = 8'b01111110; | Outputs: P=%b | Expected: P=%d",
                 1698,
                 
                 P
                 , 
                 
                 27594
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011010; B = 8'b11000010; // Expected: {'P': 5044}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011010; B = 8'b11000010; | Outputs: P=%b | Expected: P=%d",
                 1699,
                 
                 P
                 , 
                 
                 5044
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101001; B = 8'b11011011; // Expected: {'P': 8979}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101001; B = 8'b11011011; | Outputs: P=%b | Expected: P=%d",
                 1700,
                 
                 P
                 , 
                 
                 8979
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000111; B = 8'b11001010; // Expected: {'P': 27270}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000111; B = 8'b11001010; | Outputs: P=%b | Expected: P=%d",
                 1701,
                 
                 P
                 , 
                 
                 27270
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101110; B = 8'b00111100; // Expected: {'P': 6600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101110; B = 8'b00111100; | Outputs: P=%b | Expected: P=%d",
                 1702,
                 
                 P
                 , 
                 
                 6600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111010; B = 8'b01000011; // Expected: {'P': 12462}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111010; B = 8'b01000011; | Outputs: P=%b | Expected: P=%d",
                 1703,
                 
                 P
                 , 
                 
                 12462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010101; B = 8'b01001100; // Expected: {'P': 1596}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010101; B = 8'b01001100; | Outputs: P=%b | Expected: P=%d",
                 1704,
                 
                 P
                 , 
                 
                 1596
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000100; B = 8'b00010111; // Expected: {'P': 4508}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000100; B = 8'b00010111; | Outputs: P=%b | Expected: P=%d",
                 1705,
                 
                 P
                 , 
                 
                 4508
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010100; B = 8'b10001010; // Expected: {'P': 20424}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010100; B = 8'b10001010; | Outputs: P=%b | Expected: P=%d",
                 1706,
                 
                 P
                 , 
                 
                 20424
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111010; B = 8'b01000000; // Expected: {'P': 7808}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111010; B = 8'b01000000; | Outputs: P=%b | Expected: P=%d",
                 1707,
                 
                 P
                 , 
                 
                 7808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001101; B = 8'b10100100; // Expected: {'P': 2132}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001101; B = 8'b10100100; | Outputs: P=%b | Expected: P=%d",
                 1708,
                 
                 P
                 , 
                 
                 2132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010100; B = 8'b01111111; // Expected: {'P': 2540}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010100; B = 8'b01111111; | Outputs: P=%b | Expected: P=%d",
                 1709,
                 
                 P
                 , 
                 
                 2540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001101; B = 8'b11100011; // Expected: {'P': 2951}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001101; B = 8'b11100011; | Outputs: P=%b | Expected: P=%d",
                 1710,
                 
                 P
                 , 
                 
                 2951
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111000; B = 8'b10010100; // Expected: {'P': 36704}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111000; B = 8'b10010100; | Outputs: P=%b | Expected: P=%d",
                 1711,
                 
                 P
                 , 
                 
                 36704
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011110; B = 8'b00000011; // Expected: {'P': 90}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011110; B = 8'b00000011; | Outputs: P=%b | Expected: P=%d",
                 1712,
                 
                 P
                 , 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010110; B = 8'b00100011; // Expected: {'P': 3010}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010110; B = 8'b00100011; | Outputs: P=%b | Expected: P=%d",
                 1713,
                 
                 P
                 , 
                 
                 3010
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000001; B = 8'b01101111; // Expected: {'P': 111}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000001; B = 8'b01101111; | Outputs: P=%b | Expected: P=%d",
                 1714,
                 
                 P
                 , 
                 
                 111
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100001; B = 8'b10101011; // Expected: {'P': 16587}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100001; B = 8'b10101011; | Outputs: P=%b | Expected: P=%d",
                 1715,
                 
                 P
                 , 
                 
                 16587
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101010; B = 8'b01011100; // Expected: {'P': 21528}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101010; B = 8'b01011100; | Outputs: P=%b | Expected: P=%d",
                 1716,
                 
                 P
                 , 
                 
                 21528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000111; B = 8'b00011100; // Expected: {'P': 3780}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000111; B = 8'b00011100; | Outputs: P=%b | Expected: P=%d",
                 1717,
                 
                 P
                 , 
                 
                 3780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110110; B = 8'b00110000; // Expected: {'P': 2592}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110110; B = 8'b00110000; | Outputs: P=%b | Expected: P=%d",
                 1718,
                 
                 P
                 , 
                 
                 2592
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101010; B = 8'b10010111; // Expected: {'P': 6342}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101010; B = 8'b10010111; | Outputs: P=%b | Expected: P=%d",
                 1719,
                 
                 P
                 , 
                 
                 6342
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011000; B = 8'b00010010; // Expected: {'P': 3888}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011000; B = 8'b00010010; | Outputs: P=%b | Expected: P=%d",
                 1720,
                 
                 P
                 , 
                 
                 3888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111100; B = 8'b10001011; // Expected: {'P': 35028}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111100; B = 8'b10001011; | Outputs: P=%b | Expected: P=%d",
                 1721,
                 
                 P
                 , 
                 
                 35028
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001010; B = 8'b01011011; // Expected: {'P': 18382}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001010; B = 8'b01011011; | Outputs: P=%b | Expected: P=%d",
                 1722,
                 
                 P
                 , 
                 
                 18382
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101110; B = 8'b10000000; // Expected: {'P': 5888}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101110; B = 8'b10000000; | Outputs: P=%b | Expected: P=%d",
                 1723,
                 
                 P
                 , 
                 
                 5888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000010; B = 8'b11100111; // Expected: {'P': 30030}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000010; B = 8'b11100111; | Outputs: P=%b | Expected: P=%d",
                 1724,
                 
                 P
                 , 
                 
                 30030
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011001; B = 8'b01011000; // Expected: {'P': 7832}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011001; B = 8'b01011000; | Outputs: P=%b | Expected: P=%d",
                 1725,
                 
                 P
                 , 
                 
                 7832
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100101; B = 8'b11011110; // Expected: {'P': 22422}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100101; B = 8'b11011110; | Outputs: P=%b | Expected: P=%d",
                 1726,
                 
                 P
                 , 
                 
                 22422
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001100; B = 8'b11011001; // Expected: {'P': 16492}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001100; B = 8'b11011001; | Outputs: P=%b | Expected: P=%d",
                 1727,
                 
                 P
                 , 
                 
                 16492
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110011; B = 8'b11001001; // Expected: {'P': 10251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110011; B = 8'b11001001; | Outputs: P=%b | Expected: P=%d",
                 1728,
                 
                 P
                 , 
                 
                 10251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100011; B = 8'b10011110; // Expected: {'P': 35866}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100011; B = 8'b10011110; | Outputs: P=%b | Expected: P=%d",
                 1729,
                 
                 P
                 , 
                 
                 35866
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101101; B = 8'b10110011; // Expected: {'P': 19511}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101101; B = 8'b10110011; | Outputs: P=%b | Expected: P=%d",
                 1730,
                 
                 P
                 , 
                 
                 19511
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011010; B = 8'b10111111; // Expected: {'P': 17190}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011010; B = 8'b10111111; | Outputs: P=%b | Expected: P=%d",
                 1731,
                 
                 P
                 , 
                 
                 17190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011011; B = 8'b01010010; // Expected: {'P': 12710}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011011; B = 8'b01010010; | Outputs: P=%b | Expected: P=%d",
                 1732,
                 
                 P
                 , 
                 
                 12710
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010010; B = 8'b01010011; // Expected: {'P': 17430}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010010; B = 8'b01010011; | Outputs: P=%b | Expected: P=%d",
                 1733,
                 
                 P
                 , 
                 
                 17430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100000; B = 8'b10100011; // Expected: {'P': 5216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100000; B = 8'b10100011; | Outputs: P=%b | Expected: P=%d",
                 1734,
                 
                 P
                 , 
                 
                 5216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010100; B = 8'b11101011; // Expected: {'P': 4700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010100; B = 8'b11101011; | Outputs: P=%b | Expected: P=%d",
                 1735,
                 
                 P
                 , 
                 
                 4700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011100; B = 8'b11111001; // Expected: {'P': 38844}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011100; B = 8'b11111001; | Outputs: P=%b | Expected: P=%d",
                 1736,
                 
                 P
                 , 
                 
                 38844
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011111; B = 8'b00100011; // Expected: {'P': 1085}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011111; B = 8'b00100011; | Outputs: P=%b | Expected: P=%d",
                 1737,
                 
                 P
                 , 
                 
                 1085
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011111; B = 8'b11011100; // Expected: {'P': 49060}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011111; B = 8'b11011100; | Outputs: P=%b | Expected: P=%d",
                 1738,
                 
                 P
                 , 
                 
                 49060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011110; B = 8'b10100110; // Expected: {'P': 26228}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011110; B = 8'b10100110; | Outputs: P=%b | Expected: P=%d",
                 1739,
                 
                 P
                 , 
                 
                 26228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100000; B = 8'b00100101; // Expected: {'P': 3552}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100000; B = 8'b00100101; | Outputs: P=%b | Expected: P=%d",
                 1740,
                 
                 P
                 , 
                 
                 3552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101101; B = 8'b00101010; // Expected: {'P': 4578}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101101; B = 8'b00101010; | Outputs: P=%b | Expected: P=%d",
                 1741,
                 
                 P
                 , 
                 
                 4578
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000000; B = 8'b00001011; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000000; B = 8'b00001011; | Outputs: P=%b | Expected: P=%d",
                 1742,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001101; B = 8'b10110001; // Expected: {'P': 13629}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001101; B = 8'b10110001; | Outputs: P=%b | Expected: P=%d",
                 1743,
                 
                 P
                 , 
                 
                 13629
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010001; B = 8'b01001001; // Expected: {'P': 10585}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010001; B = 8'b01001001; | Outputs: P=%b | Expected: P=%d",
                 1744,
                 
                 P
                 , 
                 
                 10585
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001101; B = 8'b00010111; // Expected: {'P': 1771}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001101; B = 8'b00010111; | Outputs: P=%b | Expected: P=%d",
                 1745,
                 
                 P
                 , 
                 
                 1771
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100000; B = 8'b10110110; // Expected: {'P': 5824}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100000; B = 8'b10110110; | Outputs: P=%b | Expected: P=%d",
                 1746,
                 
                 P
                 , 
                 
                 5824
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011010; B = 8'b11110111; // Expected: {'P': 53846}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011010; B = 8'b11110111; | Outputs: P=%b | Expected: P=%d",
                 1747,
                 
                 P
                 , 
                 
                 53846
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100101; B = 8'b11011110; // Expected: {'P': 8214}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100101; B = 8'b11011110; | Outputs: P=%b | Expected: P=%d",
                 1748,
                 
                 P
                 , 
                 
                 8214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001001; B = 8'b10100100; // Expected: {'P': 1476}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001001; B = 8'b10100100; | Outputs: P=%b | Expected: P=%d",
                 1749,
                 
                 P
                 , 
                 
                 1476
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100011; B = 8'b01101001; // Expected: {'P': 23835}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100011; B = 8'b01101001; | Outputs: P=%b | Expected: P=%d",
                 1750,
                 
                 P
                 , 
                 
                 23835
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000110; B = 8'b00110110; // Expected: {'P': 10692}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000110; B = 8'b00110110; | Outputs: P=%b | Expected: P=%d",
                 1751,
                 
                 P
                 , 
                 
                 10692
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101000; B = 8'b01110101; // Expected: {'P': 27144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101000; B = 8'b01110101; | Outputs: P=%b | Expected: P=%d",
                 1752,
                 
                 P
                 , 
                 
                 27144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001111; B = 8'b01110101; // Expected: {'P': 9243}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001111; B = 8'b01110101; | Outputs: P=%b | Expected: P=%d",
                 1753,
                 
                 P
                 , 
                 
                 9243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010100; B = 8'b00010101; // Expected: {'P': 420}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010100; B = 8'b00010101; | Outputs: P=%b | Expected: P=%d",
                 1754,
                 
                 P
                 , 
                 
                 420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101110; B = 8'b11110011; // Expected: {'P': 26730}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101110; B = 8'b11110011; | Outputs: P=%b | Expected: P=%d",
                 1755,
                 
                 P
                 , 
                 
                 26730
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000111; B = 8'b10001010; // Expected: {'P': 9798}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000111; B = 8'b10001010; | Outputs: P=%b | Expected: P=%d",
                 1756,
                 
                 P
                 , 
                 
                 9798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011010; B = 8'b01011111; // Expected: {'P': 2470}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011010; B = 8'b01011111; | Outputs: P=%b | Expected: P=%d",
                 1757,
                 
                 P
                 , 
                 
                 2470
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011110; B = 8'b01101111; // Expected: {'P': 17538}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011110; B = 8'b01101111; | Outputs: P=%b | Expected: P=%d",
                 1758,
                 
                 P
                 , 
                 
                 17538
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111110; B = 8'b00000101; // Expected: {'P': 950}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111110; B = 8'b00000101; | Outputs: P=%b | Expected: P=%d",
                 1759,
                 
                 P
                 , 
                 
                 950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111100; B = 8'b00010101; // Expected: {'P': 1260}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111100; B = 8'b00010101; | Outputs: P=%b | Expected: P=%d",
                 1760,
                 
                 P
                 , 
                 
                 1260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111010; B = 8'b11110000; // Expected: {'P': 29280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111010; B = 8'b11110000; | Outputs: P=%b | Expected: P=%d",
                 1761,
                 
                 P
                 , 
                 
                 29280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100101; B = 8'b10100000; // Expected: {'P': 26400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100101; B = 8'b10100000; | Outputs: P=%b | Expected: P=%d",
                 1762,
                 
                 P
                 , 
                 
                 26400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111111; B = 8'b00000011; // Expected: {'P': 573}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111111; B = 8'b00000011; | Outputs: P=%b | Expected: P=%d",
                 1763,
                 
                 P
                 , 
                 
                 573
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010100; B = 8'b11000110; // Expected: {'P': 3960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010100; B = 8'b11000110; | Outputs: P=%b | Expected: P=%d",
                 1764,
                 
                 P
                 , 
                 
                 3960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101111; B = 8'b10001101; // Expected: {'P': 15651}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101111; B = 8'b10001101; | Outputs: P=%b | Expected: P=%d",
                 1765,
                 
                 P
                 , 
                 
                 15651
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010010; B = 8'b01000000; // Expected: {'P': 5248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010010; B = 8'b01000000; | Outputs: P=%b | Expected: P=%d",
                 1766,
                 
                 P
                 , 
                 
                 5248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111000; B = 8'b11110100; // Expected: {'P': 29280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111000; B = 8'b11110100; | Outputs: P=%b | Expected: P=%d",
                 1767,
                 
                 P
                 , 
                 
                 29280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001001; B = 8'b00011000; // Expected: {'P': 4824}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001001; B = 8'b00011000; | Outputs: P=%b | Expected: P=%d",
                 1768,
                 
                 P
                 , 
                 
                 4824
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011001; B = 8'b00101010; // Expected: {'P': 3738}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011001; B = 8'b00101010; | Outputs: P=%b | Expected: P=%d",
                 1769,
                 
                 P
                 , 
                 
                 3738
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001100; B = 8'b10000110; // Expected: {'P': 18760}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001100; B = 8'b10000110; | Outputs: P=%b | Expected: P=%d",
                 1770,
                 
                 P
                 , 
                 
                 18760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111000; B = 8'b01010011; // Expected: {'P': 20584}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111000; B = 8'b01010011; | Outputs: P=%b | Expected: P=%d",
                 1771,
                 
                 P
                 , 
                 
                 20584
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110010; B = 8'b10000001; // Expected: {'P': 6450}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110010; B = 8'b10000001; | Outputs: P=%b | Expected: P=%d",
                 1772,
                 
                 P
                 , 
                 
                 6450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100001; B = 8'b11100100; // Expected: {'P': 22116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100001; B = 8'b11100100; | Outputs: P=%b | Expected: P=%d",
                 1773,
                 
                 P
                 , 
                 
                 22116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000000; B = 8'b10100000; // Expected: {'P': 10240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000000; B = 8'b10100000; | Outputs: P=%b | Expected: P=%d",
                 1774,
                 
                 P
                 , 
                 
                 10240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010011; B = 8'b11111101; // Expected: {'P': 4807}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010011; B = 8'b11111101; | Outputs: P=%b | Expected: P=%d",
                 1775,
                 
                 P
                 , 
                 
                 4807
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110101; B = 8'b00000001; // Expected: {'P': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110101; B = 8'b00000001; | Outputs: P=%b | Expected: P=%d",
                 1776,
                 
                 P
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000100; B = 8'b01111110; // Expected: {'P': 8568}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000100; B = 8'b01111110; | Outputs: P=%b | Expected: P=%d",
                 1777,
                 
                 P
                 , 
                 
                 8568
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010001; B = 8'b11110111; // Expected: {'P': 51623}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010001; B = 8'b11110111; | Outputs: P=%b | Expected: P=%d",
                 1778,
                 
                 P
                 , 
                 
                 51623
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110000; B = 8'b00111001; // Expected: {'P': 2736}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110000; B = 8'b00111001; | Outputs: P=%b | Expected: P=%d",
                 1779,
                 
                 P
                 , 
                 
                 2736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000110; B = 8'b11011100; // Expected: {'P': 29480}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000110; B = 8'b11011100; | Outputs: P=%b | Expected: P=%d",
                 1780,
                 
                 P
                 , 
                 
                 29480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111010; B = 8'b01000100; // Expected: {'P': 3944}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111010; B = 8'b01000100; | Outputs: P=%b | Expected: P=%d",
                 1781,
                 
                 P
                 , 
                 
                 3944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101010; B = 8'b10011100; // Expected: {'P': 6552}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101010; B = 8'b10011100; | Outputs: P=%b | Expected: P=%d",
                 1782,
                 
                 P
                 , 
                 
                 6552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011110; B = 8'b10100110; // Expected: {'P': 15604}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011110; B = 8'b10100110; | Outputs: P=%b | Expected: P=%d",
                 1783,
                 
                 P
                 , 
                 
                 15604
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101010; B = 8'b10000110; // Expected: {'P': 31356}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101010; B = 8'b10000110; | Outputs: P=%b | Expected: P=%d",
                 1784,
                 
                 P
                 , 
                 
                 31356
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001010; B = 8'b10101010; // Expected: {'P': 1700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001010; B = 8'b10101010; | Outputs: P=%b | Expected: P=%d",
                 1785,
                 
                 P
                 , 
                 
                 1700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010110; B = 8'b10100111; // Expected: {'P': 35738}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010110; B = 8'b10100111; | Outputs: P=%b | Expected: P=%d",
                 1786,
                 
                 P
                 , 
                 
                 35738
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001010; B = 8'b00000110; // Expected: {'P': 828}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001010; B = 8'b00000110; | Outputs: P=%b | Expected: P=%d",
                 1787,
                 
                 P
                 , 
                 
                 828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100100; B = 8'b11100010; // Expected: {'P': 51528}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100100; B = 8'b11100010; | Outputs: P=%b | Expected: P=%d",
                 1788,
                 
                 P
                 , 
                 
                 51528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110111; B = 8'b11010000; // Expected: {'P': 11440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110111; B = 8'b11010000; | Outputs: P=%b | Expected: P=%d",
                 1789,
                 
                 P
                 , 
                 
                 11440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111011; B = 8'b00111010; // Expected: {'P': 3422}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111011; B = 8'b00111010; | Outputs: P=%b | Expected: P=%d",
                 1790,
                 
                 P
                 , 
                 
                 3422
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110111; B = 8'b10100110; // Expected: {'P': 30378}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110111; B = 8'b10100110; | Outputs: P=%b | Expected: P=%d",
                 1791,
                 
                 P
                 , 
                 
                 30378
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001101; B = 8'b01011010; // Expected: {'P': 12690}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001101; B = 8'b01011010; | Outputs: P=%b | Expected: P=%d",
                 1792,
                 
                 P
                 , 
                 
                 12690
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010111; B = 8'b10111111; // Expected: {'P': 16617}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010111; B = 8'b10111111; | Outputs: P=%b | Expected: P=%d",
                 1793,
                 
                 P
                 , 
                 
                 16617
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111111; B = 8'b11100111; // Expected: {'P': 44121}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111111; B = 8'b11100111; | Outputs: P=%b | Expected: P=%d",
                 1794,
                 
                 P
                 , 
                 
                 44121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000001; B = 8'b11111110; // Expected: {'P': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000001; B = 8'b11111110; | Outputs: P=%b | Expected: P=%d",
                 1795,
                 
                 P
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110101; B = 8'b11010010; // Expected: {'P': 11130}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110101; B = 8'b11010010; | Outputs: P=%b | Expected: P=%d",
                 1796,
                 
                 P
                 , 
                 
                 11130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000110; B = 8'b01010100; // Expected: {'P': 16632}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000110; B = 8'b01010100; | Outputs: P=%b | Expected: P=%d",
                 1797,
                 
                 P
                 , 
                 
                 16632
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011011; B = 8'b00011010; // Expected: {'P': 5694}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011011; B = 8'b00011010; | Outputs: P=%b | Expected: P=%d",
                 1798,
                 
                 P
                 , 
                 
                 5694
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101100; B = 8'b00101110; // Expected: {'P': 7912}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101100; B = 8'b00101110; | Outputs: P=%b | Expected: P=%d",
                 1799,
                 
                 P
                 , 
                 
                 7912
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101011; B = 8'b01110011; // Expected: {'P': 19665}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101011; B = 8'b01110011; | Outputs: P=%b | Expected: P=%d",
                 1800,
                 
                 P
                 , 
                 
                 19665
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010101; B = 8'b00101101; // Expected: {'P': 9585}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010101; B = 8'b00101101; | Outputs: P=%b | Expected: P=%d",
                 1801,
                 
                 P
                 , 
                 
                 9585
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011010; B = 8'b01010101; // Expected: {'P': 13090}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011010; B = 8'b01010101; | Outputs: P=%b | Expected: P=%d",
                 1802,
                 
                 P
                 , 
                 
                 13090
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100001; B = 8'b01110111; // Expected: {'P': 19159}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100001; B = 8'b01110111; | Outputs: P=%b | Expected: P=%d",
                 1803,
                 
                 P
                 , 
                 
                 19159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011111; B = 8'b00111011; // Expected: {'P': 9381}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011111; B = 8'b00111011; | Outputs: P=%b | Expected: P=%d",
                 1804,
                 
                 P
                 , 
                 
                 9381
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001011; B = 8'b01010011; // Expected: {'P': 913}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001011; B = 8'b01010011; | Outputs: P=%b | Expected: P=%d",
                 1805,
                 
                 P
                 , 
                 
                 913
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101010; B = 8'b01010011; // Expected: {'P': 3486}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101010; B = 8'b01010011; | Outputs: P=%b | Expected: P=%d",
                 1806,
                 
                 P
                 , 
                 
                 3486
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000101; B = 8'b00010001; // Expected: {'P': 3349}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000101; B = 8'b00010001; | Outputs: P=%b | Expected: P=%d",
                 1807,
                 
                 P
                 , 
                 
                 3349
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011011; B = 8'b11011100; // Expected: {'P': 34100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011011; B = 8'b11011100; | Outputs: P=%b | Expected: P=%d",
                 1808,
                 
                 P
                 , 
                 
                 34100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010111; B = 8'b00100101; // Expected: {'P': 851}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010111; B = 8'b00100101; | Outputs: P=%b | Expected: P=%d",
                 1809,
                 
                 P
                 , 
                 
                 851
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111001; B = 8'b10110001; // Expected: {'P': 44073}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111001; B = 8'b10110001; | Outputs: P=%b | Expected: P=%d",
                 1810,
                 
                 P
                 , 
                 
                 44073
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000001; B = 8'b01111011; // Expected: {'P': 123}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000001; B = 8'b01111011; | Outputs: P=%b | Expected: P=%d",
                 1811,
                 
                 P
                 , 
                 
                 123
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110111; B = 8'b11101101; // Expected: {'P': 58539}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110111; B = 8'b11101101; | Outputs: P=%b | Expected: P=%d",
                 1812,
                 
                 P
                 , 
                 
                 58539
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000101; B = 8'b01110011; // Expected: {'P': 15295}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000101; B = 8'b01110011; | Outputs: P=%b | Expected: P=%d",
                 1813,
                 
                 P
                 , 
                 
                 15295
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101001; B = 8'b11011111; // Expected: {'P': 37687}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101001; B = 8'b11011111; | Outputs: P=%b | Expected: P=%d",
                 1814,
                 
                 P
                 , 
                 
                 37687
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010011; B = 8'b01011000; // Expected: {'P': 1672}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010011; B = 8'b01011000; | Outputs: P=%b | Expected: P=%d",
                 1815,
                 
                 P
                 , 
                 
                 1672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110010; B = 8'b01100110; // Expected: {'P': 24684}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110010; B = 8'b01100110; | Outputs: P=%b | Expected: P=%d",
                 1816,
                 
                 P
                 , 
                 
                 24684
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100110; B = 8'b00010100; // Expected: {'P': 760}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100110; B = 8'b00010100; | Outputs: P=%b | Expected: P=%d",
                 1817,
                 
                 P
                 , 
                 
                 760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011101; B = 8'b00111100; // Expected: {'P': 5580}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011101; B = 8'b00111100; | Outputs: P=%b | Expected: P=%d",
                 1818,
                 
                 P
                 , 
                 
                 5580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011101; B = 8'b11101100; // Expected: {'P': 37052}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011101; B = 8'b11101100; | Outputs: P=%b | Expected: P=%d",
                 1819,
                 
                 P
                 , 
                 
                 37052
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011010; B = 8'b11100011; // Expected: {'P': 20430}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011010; B = 8'b11100011; | Outputs: P=%b | Expected: P=%d",
                 1820,
                 
                 P
                 , 
                 
                 20430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111000; B = 8'b10111111; // Expected: {'P': 22920}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111000; B = 8'b10111111; | Outputs: P=%b | Expected: P=%d",
                 1821,
                 
                 P
                 , 
                 
                 22920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100000; B = 8'b10000010; // Expected: {'P': 20800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100000; B = 8'b10000010; | Outputs: P=%b | Expected: P=%d",
                 1822,
                 
                 P
                 , 
                 
                 20800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001011; B = 8'b00110010; // Expected: {'P': 10150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001011; B = 8'b00110010; | Outputs: P=%b | Expected: P=%d",
                 1823,
                 
                 P
                 , 
                 
                 10150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011001; B = 8'b00111100; // Expected: {'P': 5340}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011001; B = 8'b00111100; | Outputs: P=%b | Expected: P=%d",
                 1824,
                 
                 P
                 , 
                 
                 5340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000101; B = 8'b00101001; // Expected: {'P': 5453}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000101; B = 8'b00101001; | Outputs: P=%b | Expected: P=%d",
                 1825,
                 
                 P
                 , 
                 
                 5453
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011000; B = 8'b01010011; // Expected: {'P': 12616}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011000; B = 8'b01010011; | Outputs: P=%b | Expected: P=%d",
                 1826,
                 
                 P
                 , 
                 
                 12616
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010101; B = 8'b00010010; // Expected: {'P': 378}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010101; B = 8'b00010010; | Outputs: P=%b | Expected: P=%d",
                 1827,
                 
                 P
                 , 
                 
                 378
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100100; B = 8'b11111101; // Expected: {'P': 57684}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100100; B = 8'b11111101; | Outputs: P=%b | Expected: P=%d",
                 1828,
                 
                 P
                 , 
                 
                 57684
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010011; B = 8'b00000011; // Expected: {'P': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010011; B = 8'b00000011; | Outputs: P=%b | Expected: P=%d",
                 1829,
                 
                 P
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011100; B = 8'b00000110; // Expected: {'P': 168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011100; B = 8'b00000110; | Outputs: P=%b | Expected: P=%d",
                 1830,
                 
                 P
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010001; B = 8'b01000011; // Expected: {'P': 9715}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010001; B = 8'b01000011; | Outputs: P=%b | Expected: P=%d",
                 1831,
                 
                 P
                 , 
                 
                 9715
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000001; B = 8'b01010110; // Expected: {'P': 16598}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000001; B = 8'b01010110; | Outputs: P=%b | Expected: P=%d",
                 1832,
                 
                 P
                 , 
                 
                 16598
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000011; B = 8'b01101100; // Expected: {'P': 21060}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000011; B = 8'b01101100; | Outputs: P=%b | Expected: P=%d",
                 1833,
                 
                 P
                 , 
                 
                 21060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000111; B = 8'b01101001; // Expected: {'P': 20895}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000111; B = 8'b01101001; | Outputs: P=%b | Expected: P=%d",
                 1834,
                 
                 P
                 , 
                 
                 20895
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010101; B = 8'b10011011; // Expected: {'P': 33015}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010101; B = 8'b10011011; | Outputs: P=%b | Expected: P=%d",
                 1835,
                 
                 P
                 , 
                 
                 33015
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101010; B = 8'b00101111; // Expected: {'P': 7990}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101010; B = 8'b00101111; | Outputs: P=%b | Expected: P=%d",
                 1836,
                 
                 P
                 , 
                 
                 7990
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100001; B = 8'b00110111; // Expected: {'P': 8855}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100001; B = 8'b00110111; | Outputs: P=%b | Expected: P=%d",
                 1837,
                 
                 P
                 , 
                 
                 8855
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110101; B = 8'b01000110; // Expected: {'P': 8190}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110101; B = 8'b01000110; | Outputs: P=%b | Expected: P=%d",
                 1838,
                 
                 P
                 , 
                 
                 8190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000010; B = 8'b11101100; // Expected: {'P': 30680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000010; B = 8'b11101100; | Outputs: P=%b | Expected: P=%d",
                 1839,
                 
                 P
                 , 
                 
                 30680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010011; B = 8'b00001111; // Expected: {'P': 2205}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010011; B = 8'b00001111; | Outputs: P=%b | Expected: P=%d",
                 1840,
                 
                 P
                 , 
                 
                 2205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010000; B = 8'b00110100; // Expected: {'P': 832}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010000; B = 8'b00110100; | Outputs: P=%b | Expected: P=%d",
                 1841,
                 
                 P
                 , 
                 
                 832
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011110; B = 8'b11001101; // Expected: {'P': 32390}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011110; B = 8'b11001101; | Outputs: P=%b | Expected: P=%d",
                 1842,
                 
                 P
                 , 
                 
                 32390
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111101; B = 8'b01011111; // Expected: {'P': 17955}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111101; B = 8'b01011111; | Outputs: P=%b | Expected: P=%d",
                 1843,
                 
                 P
                 , 
                 
                 17955
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111100; B = 8'b01000110; // Expected: {'P': 4200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111100; B = 8'b01000110; | Outputs: P=%b | Expected: P=%d",
                 1844,
                 
                 P
                 , 
                 
                 4200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010010; B = 8'b00000110; // Expected: {'P': 492}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010010; B = 8'b00000110; | Outputs: P=%b | Expected: P=%d",
                 1845,
                 
                 P
                 , 
                 
                 492
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111011; B = 8'b11001010; // Expected: {'P': 24846}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111011; B = 8'b11001010; | Outputs: P=%b | Expected: P=%d",
                 1846,
                 
                 P
                 , 
                 
                 24846
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000111; B = 8'b11110001; // Expected: {'P': 1687}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000111; B = 8'b11110001; | Outputs: P=%b | Expected: P=%d",
                 1847,
                 
                 P
                 , 
                 
                 1687
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000001; B = 8'b01011101; // Expected: {'P': 6045}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000001; B = 8'b01011101; | Outputs: P=%b | Expected: P=%d",
                 1848,
                 
                 P
                 , 
                 
                 6045
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010000; B = 8'b01001101; // Expected: {'P': 16016}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010000; B = 8'b01001101; | Outputs: P=%b | Expected: P=%d",
                 1849,
                 
                 P
                 , 
                 
                 16016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011000; B = 8'b11101110; // Expected: {'P': 5712}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011000; B = 8'b11101110; | Outputs: P=%b | Expected: P=%d",
                 1850,
                 
                 P
                 , 
                 
                 5712
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010100; B = 8'b00110111; // Expected: {'P': 8140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010100; B = 8'b00110111; | Outputs: P=%b | Expected: P=%d",
                 1851,
                 
                 P
                 , 
                 
                 8140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111011; B = 8'b11100111; // Expected: {'P': 43197}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111011; B = 8'b11100111; | Outputs: P=%b | Expected: P=%d",
                 1852,
                 
                 P
                 , 
                 
                 43197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010010; B = 8'b11111100; // Expected: {'P': 52920}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010010; B = 8'b11111100; | Outputs: P=%b | Expected: P=%d",
                 1853,
                 
                 P
                 , 
                 
                 52920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101111; B = 8'b01010111; // Expected: {'P': 15225}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101111; B = 8'b01010111; | Outputs: P=%b | Expected: P=%d",
                 1854,
                 
                 P
                 , 
                 
                 15225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010001; B = 8'b11000011; // Expected: {'P': 3315}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010001; B = 8'b11000011; | Outputs: P=%b | Expected: P=%d",
                 1855,
                 
                 P
                 , 
                 
                 3315
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110000; B = 8'b11001001; // Expected: {'P': 9648}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110000; B = 8'b11001001; | Outputs: P=%b | Expected: P=%d",
                 1856,
                 
                 P
                 , 
                 
                 9648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000000; B = 8'b11100110; // Expected: {'P': 44160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000000; B = 8'b11100110; | Outputs: P=%b | Expected: P=%d",
                 1857,
                 
                 P
                 , 
                 
                 44160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000111; B = 8'b10100110; // Expected: {'P': 11786}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000111; B = 8'b10100110; | Outputs: P=%b | Expected: P=%d",
                 1858,
                 
                 P
                 , 
                 
                 11786
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101010; B = 8'b10101001; // Expected: {'P': 7098}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101010; B = 8'b10101001; | Outputs: P=%b | Expected: P=%d",
                 1859,
                 
                 P
                 , 
                 
                 7098
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011100; B = 8'b10001001; // Expected: {'P': 21372}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011100; B = 8'b10001001; | Outputs: P=%b | Expected: P=%d",
                 1860,
                 
                 P
                 , 
                 
                 21372
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010101; B = 8'b01101111; // Expected: {'P': 2331}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010101; B = 8'b01101111; | Outputs: P=%b | Expected: P=%d",
                 1861,
                 
                 P
                 , 
                 
                 2331
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011010; B = 8'b11001111; // Expected: {'P': 45126}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011010; B = 8'b11001111; | Outputs: P=%b | Expected: P=%d",
                 1862,
                 
                 P
                 , 
                 
                 45126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111111; B = 8'b11000001; // Expected: {'P': 12159}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111111; B = 8'b11000001; | Outputs: P=%b | Expected: P=%d",
                 1863,
                 
                 P
                 , 
                 
                 12159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001110; B = 8'b00011011; // Expected: {'P': 3834}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001110; B = 8'b00011011; | Outputs: P=%b | Expected: P=%d",
                 1864,
                 
                 P
                 , 
                 
                 3834
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100000; B = 8'b10011000; // Expected: {'P': 24320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100000; B = 8'b10011000; | Outputs: P=%b | Expected: P=%d",
                 1865,
                 
                 P
                 , 
                 
                 24320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101110; B = 8'b00001000; // Expected: {'P': 1392}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101110; B = 8'b00001000; | Outputs: P=%b | Expected: P=%d",
                 1866,
                 
                 P
                 , 
                 
                 1392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110011; B = 8'b11001110; // Expected: {'P': 10506}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110011; B = 8'b11001110; | Outputs: P=%b | Expected: P=%d",
                 1867,
                 
                 P
                 , 
                 
                 10506
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000011; B = 8'b11001100; // Expected: {'P': 26724}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000011; B = 8'b11001100; | Outputs: P=%b | Expected: P=%d",
                 1868,
                 
                 P
                 , 
                 
                 26724
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000010; B = 8'b00010100; // Expected: {'P': 2600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000010; B = 8'b00010100; | Outputs: P=%b | Expected: P=%d",
                 1869,
                 
                 P
                 , 
                 
                 2600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110101; B = 8'b00001101; // Expected: {'P': 1521}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110101; B = 8'b00001101; | Outputs: P=%b | Expected: P=%d",
                 1870,
                 
                 P
                 , 
                 
                 1521
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100111; B = 8'b00100001; // Expected: {'P': 1287}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100111; B = 8'b00100001; | Outputs: P=%b | Expected: P=%d",
                 1871,
                 
                 P
                 , 
                 
                 1287
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001101; B = 8'b01000101; // Expected: {'P': 5313}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001101; B = 8'b01000101; | Outputs: P=%b | Expected: P=%d",
                 1872,
                 
                 P
                 , 
                 
                 5313
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001101; B = 8'b10001000; // Expected: {'P': 27880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001101; B = 8'b10001000; | Outputs: P=%b | Expected: P=%d",
                 1873,
                 
                 P
                 , 
                 
                 27880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101100; B = 8'b11101011; // Expected: {'P': 40420}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101100; B = 8'b11101011; | Outputs: P=%b | Expected: P=%d",
                 1874,
                 
                 P
                 , 
                 
                 40420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000001; B = 8'b00110111; // Expected: {'P': 3575}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000001; B = 8'b00110111; | Outputs: P=%b | Expected: P=%d",
                 1875,
                 
                 P
                 , 
                 
                 3575
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100001; B = 8'b11101000; // Expected: {'P': 22504}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100001; B = 8'b11101000; | Outputs: P=%b | Expected: P=%d",
                 1876,
                 
                 P
                 , 
                 
                 22504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110100; B = 8'b00011111; // Expected: {'P': 5580}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110100; B = 8'b00011111; | Outputs: P=%b | Expected: P=%d",
                 1877,
                 
                 P
                 , 
                 
                 5580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010010; B = 8'b01110110; // Expected: {'P': 9676}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010010; B = 8'b01110110; | Outputs: P=%b | Expected: P=%d",
                 1878,
                 
                 P
                 , 
                 
                 9676
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001011; B = 8'b11110001; // Expected: {'P': 2651}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001011; B = 8'b11110001; | Outputs: P=%b | Expected: P=%d",
                 1879,
                 
                 P
                 , 
                 
                 2651
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111000; B = 8'b10110011; // Expected: {'P': 44392}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111000; B = 8'b10110011; | Outputs: P=%b | Expected: P=%d",
                 1880,
                 
                 P
                 , 
                 
                 44392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101101; B = 8'b00100100; // Expected: {'P': 6228}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101101; B = 8'b00100100; | Outputs: P=%b | Expected: P=%d",
                 1881,
                 
                 P
                 , 
                 
                 6228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110000; B = 8'b10111100; // Expected: {'P': 33088}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110000; B = 8'b10111100; | Outputs: P=%b | Expected: P=%d",
                 1882,
                 
                 P
                 , 
                 
                 33088
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011011; B = 8'b00001010; // Expected: {'P': 2190}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011011; B = 8'b00001010; | Outputs: P=%b | Expected: P=%d",
                 1883,
                 
                 P
                 , 
                 
                 2190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001110; B = 8'b10011110; // Expected: {'P': 22436}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001110; B = 8'b10011110; | Outputs: P=%b | Expected: P=%d",
                 1884,
                 
                 P
                 , 
                 
                 22436
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010111; B = 8'b11001001; // Expected: {'P': 43215}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010111; B = 8'b11001001; | Outputs: P=%b | Expected: P=%d",
                 1885,
                 
                 P
                 , 
                 
                 43215
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110111; B = 8'b00101111; // Expected: {'P': 11609}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110111; B = 8'b00101111; | Outputs: P=%b | Expected: P=%d",
                 1886,
                 
                 P
                 , 
                 
                 11609
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100110; B = 8'b11110100; // Expected: {'P': 40504}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100110; B = 8'b11110100; | Outputs: P=%b | Expected: P=%d",
                 1887,
                 
                 P
                 , 
                 
                 40504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000110; B = 8'b00100100; // Expected: {'P': 7128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000110; B = 8'b00100100; | Outputs: P=%b | Expected: P=%d",
                 1888,
                 
                 P
                 , 
                 
                 7128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101000; B = 8'b00000101; // Expected: {'P': 840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101000; B = 8'b00000101; | Outputs: P=%b | Expected: P=%d",
                 1889,
                 
                 P
                 , 
                 
                 840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100101; B = 8'b01100010; // Expected: {'P': 22442}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100101; B = 8'b01100010; | Outputs: P=%b | Expected: P=%d",
                 1890,
                 
                 P
                 , 
                 
                 22442
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001101; B = 8'b11001011; // Expected: {'P': 15631}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001101; B = 8'b11001011; | Outputs: P=%b | Expected: P=%d",
                 1891,
                 
                 P
                 , 
                 
                 15631
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011100; B = 8'b00011011; // Expected: {'P': 5940}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011100; B = 8'b00011011; | Outputs: P=%b | Expected: P=%d",
                 1892,
                 
                 P
                 , 
                 
                 5940
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100001; B = 8'b11110001; // Expected: {'P': 54225}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100001; B = 8'b11110001; | Outputs: P=%b | Expected: P=%d",
                 1893,
                 
                 P
                 , 
                 
                 54225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111010; B = 8'b00100110; // Expected: {'P': 4636}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111010; B = 8'b00100110; | Outputs: P=%b | Expected: P=%d",
                 1894,
                 
                 P
                 , 
                 
                 4636
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101000; B = 8'b11100001; // Expected: {'P': 23400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101000; B = 8'b11100001; | Outputs: P=%b | Expected: P=%d",
                 1895,
                 
                 P
                 , 
                 
                 23400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001101; B = 8'b11101111; // Expected: {'P': 18403}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001101; B = 8'b11101111; | Outputs: P=%b | Expected: P=%d",
                 1896,
                 
                 P
                 , 
                 
                 18403
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001011; B = 8'b01110000; // Expected: {'P': 1232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001011; B = 8'b01110000; | Outputs: P=%b | Expected: P=%d",
                 1897,
                 
                 P
                 , 
                 
                 1232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000010; B = 8'b10101010; // Expected: {'P': 340}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000010; B = 8'b10101010; | Outputs: P=%b | Expected: P=%d",
                 1898,
                 
                 P
                 , 
                 
                 340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010000; B = 8'b11110011; // Expected: {'P': 3888}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010000; B = 8'b11110011; | Outputs: P=%b | Expected: P=%d",
                 1899,
                 
                 P
                 , 
                 
                 3888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101110; B = 8'b01111100; // Expected: {'P': 21576}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101110; B = 8'b01111100; | Outputs: P=%b | Expected: P=%d",
                 1900,
                 
                 P
                 , 
                 
                 21576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110001; B = 8'b00101100; // Expected: {'P': 2156}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110001; B = 8'b00101100; | Outputs: P=%b | Expected: P=%d",
                 1901,
                 
                 P
                 , 
                 
                 2156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000000; B = 8'b11011010; // Expected: {'P': 13952}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000000; B = 8'b11011010; | Outputs: P=%b | Expected: P=%d",
                 1902,
                 
                 P
                 , 
                 
                 13952
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101100; B = 8'b11001110; // Expected: {'P': 22248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101100; B = 8'b11001110; | Outputs: P=%b | Expected: P=%d",
                 1903,
                 
                 P
                 , 
                 
                 22248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001111; B = 8'b00010100; // Expected: {'P': 2860}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001111; B = 8'b00010100; | Outputs: P=%b | Expected: P=%d",
                 1904,
                 
                 P
                 , 
                 
                 2860
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001010; B = 8'b11001110; // Expected: {'P': 2060}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001010; B = 8'b11001110; | Outputs: P=%b | Expected: P=%d",
                 1905,
                 
                 P
                 , 
                 
                 2060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000001; B = 8'b00001010; // Expected: {'P': 650}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000001; B = 8'b00001010; | Outputs: P=%b | Expected: P=%d",
                 1906,
                 
                 P
                 , 
                 
                 650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011001; B = 8'b01001001; // Expected: {'P': 6497}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011001; B = 8'b01001001; | Outputs: P=%b | Expected: P=%d",
                 1907,
                 
                 P
                 , 
                 
                 6497
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110010; B = 8'b11000011; // Expected: {'P': 22230}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110010; B = 8'b11000011; | Outputs: P=%b | Expected: P=%d",
                 1908,
                 
                 P
                 , 
                 
                 22230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001000; B = 8'b10011111; // Expected: {'P': 1272}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001000; B = 8'b10011111; | Outputs: P=%b | Expected: P=%d",
                 1909,
                 
                 P
                 , 
                 
                 1272
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110110; B = 8'b00101000; // Expected: {'P': 2160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110110; B = 8'b00101000; | Outputs: P=%b | Expected: P=%d",
                 1910,
                 
                 P
                 , 
                 
                 2160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101111; B = 8'b00100001; // Expected: {'P': 5775}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101111; B = 8'b00100001; | Outputs: P=%b | Expected: P=%d",
                 1911,
                 
                 P
                 , 
                 
                 5775
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100100; B = 8'b01101111; // Expected: {'P': 25308}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100100; B = 8'b01101111; | Outputs: P=%b | Expected: P=%d",
                 1912,
                 
                 P
                 , 
                 
                 25308
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000111; B = 8'b01000111; // Expected: {'P': 5041}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000111; B = 8'b01000111; | Outputs: P=%b | Expected: P=%d",
                 1913,
                 
                 P
                 , 
                 
                 5041
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001100; B = 8'b00110101; // Expected: {'P': 7420}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001100; B = 8'b00110101; | Outputs: P=%b | Expected: P=%d",
                 1914,
                 
                 P
                 , 
                 
                 7420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110100; B = 8'b11001110; // Expected: {'P': 10712}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110100; B = 8'b11001110; | Outputs: P=%b | Expected: P=%d",
                 1915,
                 
                 P
                 , 
                 
                 10712
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110010; B = 8'b10001111; // Expected: {'P': 16302}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110010; B = 8'b10001111; | Outputs: P=%b | Expected: P=%d",
                 1916,
                 
                 P
                 , 
                 
                 16302
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101101; B = 8'b11111110; // Expected: {'P': 27686}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101101; B = 8'b11111110; | Outputs: P=%b | Expected: P=%d",
                 1917,
                 
                 P
                 , 
                 
                 27686
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110010; B = 8'b11010010; // Expected: {'P': 10500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110010; B = 8'b11010010; | Outputs: P=%b | Expected: P=%d",
                 1918,
                 
                 P
                 , 
                 
                 10500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101111; B = 8'b01110100; // Expected: {'P': 12876}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101111; B = 8'b01110100; | Outputs: P=%b | Expected: P=%d",
                 1919,
                 
                 P
                 , 
                 
                 12876
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001110; B = 8'b01110000; // Expected: {'P': 8736}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001110; B = 8'b01110000; | Outputs: P=%b | Expected: P=%d",
                 1920,
                 
                 P
                 , 
                 
                 8736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110001; B = 8'b01000000; // Expected: {'P': 7232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110001; B = 8'b01000000; | Outputs: P=%b | Expected: P=%d",
                 1921,
                 
                 P
                 , 
                 
                 7232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011110; B = 8'b10101000; // Expected: {'P': 5040}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011110; B = 8'b10101000; | Outputs: P=%b | Expected: P=%d",
                 1922,
                 
                 P
                 , 
                 
                 5040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101110; B = 8'b10110010; // Expected: {'P': 8188}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101110; B = 8'b10110010; | Outputs: P=%b | Expected: P=%d",
                 1923,
                 
                 P
                 , 
                 
                 8188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110110; B = 8'b01101111; // Expected: {'P': 27306}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110110; B = 8'b01101111; | Outputs: P=%b | Expected: P=%d",
                 1924,
                 
                 P
                 , 
                 
                 27306
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001111; B = 8'b00101011; // Expected: {'P': 6149}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001111; B = 8'b00101011; | Outputs: P=%b | Expected: P=%d",
                 1925,
                 
                 P
                 , 
                 
                 6149
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001010; B = 8'b00110000; // Expected: {'P': 6624}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001010; B = 8'b00110000; | Outputs: P=%b | Expected: P=%d",
                 1926,
                 
                 P
                 , 
                 
                 6624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101111; B = 8'b11101101; // Expected: {'P': 11139}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101111; B = 8'b11101101; | Outputs: P=%b | Expected: P=%d",
                 1927,
                 
                 P
                 , 
                 
                 11139
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010011; B = 8'b10000011; // Expected: {'P': 19257}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010011; B = 8'b10000011; | Outputs: P=%b | Expected: P=%d",
                 1928,
                 
                 P
                 , 
                 
                 19257
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110111; B = 8'b01110110; // Expected: {'P': 21594}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110111; B = 8'b01110110; | Outputs: P=%b | Expected: P=%d",
                 1929,
                 
                 P
                 , 
                 
                 21594
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110011; B = 8'b01110100; // Expected: {'P': 28188}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110011; B = 8'b01110100; | Outputs: P=%b | Expected: P=%d",
                 1930,
                 
                 P
                 , 
                 
                 28188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101001; B = 8'b10011110; // Expected: {'P': 16590}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101001; B = 8'b10011110; | Outputs: P=%b | Expected: P=%d",
                 1931,
                 
                 P
                 , 
                 
                 16590
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010010; B = 8'b10101001; // Expected: {'P': 35490}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010010; B = 8'b10101001; | Outputs: P=%b | Expected: P=%d",
                 1932,
                 
                 P
                 , 
                 
                 35490
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101100; B = 8'b11111011; // Expected: {'P': 59236}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101100; B = 8'b11111011; | Outputs: P=%b | Expected: P=%d",
                 1933,
                 
                 P
                 , 
                 
                 59236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101110; B = 8'b10101110; // Expected: {'P': 41412}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101110; B = 8'b10101110; | Outputs: P=%b | Expected: P=%d",
                 1934,
                 
                 P
                 , 
                 
                 41412
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111001; B = 8'b01100010; // Expected: {'P': 5586}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111001; B = 8'b01100010; | Outputs: P=%b | Expected: P=%d",
                 1935,
                 
                 P
                 , 
                 
                 5586
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111000; B = 8'b11110111; // Expected: {'P': 61256}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111000; B = 8'b11110111; | Outputs: P=%b | Expected: P=%d",
                 1936,
                 
                 P
                 , 
                 
                 61256
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001011; B = 8'b10110000; // Expected: {'P': 1936}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001011; B = 8'b10110000; | Outputs: P=%b | Expected: P=%d",
                 1937,
                 
                 P
                 , 
                 
                 1936
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101001; B = 8'b01111010; // Expected: {'P': 28426}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101001; B = 8'b01111010; | Outputs: P=%b | Expected: P=%d",
                 1938,
                 
                 P
                 , 
                 
                 28426
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011010; B = 8'b11110101; // Expected: {'P': 53410}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011010; B = 8'b11110101; | Outputs: P=%b | Expected: P=%d",
                 1939,
                 
                 P
                 , 
                 
                 53410
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011101; B = 8'b01000011; // Expected: {'P': 6231}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011101; B = 8'b01000011; | Outputs: P=%b | Expected: P=%d",
                 1940,
                 
                 P
                 , 
                 
                 6231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010101; B = 8'b00001011; // Expected: {'P': 1639}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010101; B = 8'b00001011; | Outputs: P=%b | Expected: P=%d",
                 1941,
                 
                 P
                 , 
                 
                 1639
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100111; B = 8'b11111100; // Expected: {'P': 9828}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100111; B = 8'b11111100; | Outputs: P=%b | Expected: P=%d",
                 1942,
                 
                 P
                 , 
                 
                 9828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001100; B = 8'b11001110; // Expected: {'P': 15656}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001100; B = 8'b11001110; | Outputs: P=%b | Expected: P=%d",
                 1943,
                 
                 P
                 , 
                 
                 15656
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000100; B = 8'b01100100; // Expected: {'P': 400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000100; B = 8'b01100100; | Outputs: P=%b | Expected: P=%d",
                 1944,
                 
                 P
                 , 
                 
                 400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100011; B = 8'b01011101; // Expected: {'P': 15159}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100011; B = 8'b01011101; | Outputs: P=%b | Expected: P=%d",
                 1945,
                 
                 P
                 , 
                 
                 15159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101101; B = 8'b11000000; // Expected: {'P': 33216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101101; B = 8'b11000000; | Outputs: P=%b | Expected: P=%d",
                 1946,
                 
                 P
                 , 
                 
                 33216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111101; B = 8'b00010110; // Expected: {'P': 5566}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111101; B = 8'b00010110; | Outputs: P=%b | Expected: P=%d",
                 1947,
                 
                 P
                 , 
                 
                 5566
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100001; B = 8'b00010000; // Expected: {'P': 1552}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100001; B = 8'b00010000; | Outputs: P=%b | Expected: P=%d",
                 1948,
                 
                 P
                 , 
                 
                 1552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101000; B = 8'b11000011; // Expected: {'P': 32760}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101000; B = 8'b11000011; | Outputs: P=%b | Expected: P=%d",
                 1949,
                 
                 P
                 , 
                 
                 32760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101011; B = 8'b00110011; // Expected: {'P': 2193}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101011; B = 8'b00110011; | Outputs: P=%b | Expected: P=%d",
                 1950,
                 
                 P
                 , 
                 
                 2193
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001100; B = 8'b00011110; // Expected: {'P': 4200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001100; B = 8'b00011110; | Outputs: P=%b | Expected: P=%d",
                 1951,
                 
                 P
                 , 
                 
                 4200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011010; B = 8'b11000001; // Expected: {'P': 29722}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011010; B = 8'b11000001; | Outputs: P=%b | Expected: P=%d",
                 1952,
                 
                 P
                 , 
                 
                 29722
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100111; B = 8'b11001000; // Expected: {'P': 20600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100111; B = 8'b11001000; | Outputs: P=%b | Expected: P=%d",
                 1953,
                 
                 P
                 , 
                 
                 20600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100010; B = 8'b11000100; // Expected: {'P': 44296}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100010; B = 8'b11000100; | Outputs: P=%b | Expected: P=%d",
                 1954,
                 
                 P
                 , 
                 
                 44296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011000; B = 8'b10011101; // Expected: {'P': 33912}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011000; B = 8'b10011101; | Outputs: P=%b | Expected: P=%d",
                 1955,
                 
                 P
                 , 
                 
                 33912
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100000; B = 8'b11110101; // Expected: {'P': 23520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100000; B = 8'b11110101; | Outputs: P=%b | Expected: P=%d",
                 1956,
                 
                 P
                 , 
                 
                 23520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100010; B = 8'b00101101; // Expected: {'P': 4410}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100010; B = 8'b00101101; | Outputs: P=%b | Expected: P=%d",
                 1957,
                 
                 P
                 , 
                 
                 4410
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101111; B = 8'b10010101; // Expected: {'P': 16539}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101111; B = 8'b10010101; | Outputs: P=%b | Expected: P=%d",
                 1958,
                 
                 P
                 , 
                 
                 16539
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101011; B = 8'b01100110; // Expected: {'P': 23970}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101011; B = 8'b01100110; | Outputs: P=%b | Expected: P=%d",
                 1959,
                 
                 P
                 , 
                 
                 23970
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001000; B = 8'b00001000; // Expected: {'P': 1600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001000; B = 8'b00001000; | Outputs: P=%b | Expected: P=%d",
                 1960,
                 
                 P
                 , 
                 
                 1600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111110; B = 8'b11101100; // Expected: {'P': 14632}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111110; B = 8'b11101100; | Outputs: P=%b | Expected: P=%d",
                 1961,
                 
                 P
                 , 
                 
                 14632
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001010; B = 8'b11111111; // Expected: {'P': 51510}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001010; B = 8'b11111111; | Outputs: P=%b | Expected: P=%d",
                 1962,
                 
                 P
                 , 
                 
                 51510
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010111; B = 8'b01100111; // Expected: {'P': 15553}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010111; B = 8'b01100111; | Outputs: P=%b | Expected: P=%d",
                 1963,
                 
                 P
                 , 
                 
                 15553
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001000; B = 8'b11101110; // Expected: {'P': 32368}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001000; B = 8'b11101110; | Outputs: P=%b | Expected: P=%d",
                 1964,
                 
                 P
                 , 
                 
                 32368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000001; B = 8'b10110101; // Expected: {'P': 181}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000001; B = 8'b10110101; | Outputs: P=%b | Expected: P=%d",
                 1965,
                 
                 P
                 , 
                 
                 181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010101; B = 8'b00100111; // Expected: {'P': 8307}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010101; B = 8'b00100111; | Outputs: P=%b | Expected: P=%d",
                 1966,
                 
                 P
                 , 
                 
                 8307
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010001; B = 8'b01100100; // Expected: {'P': 20900}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010001; B = 8'b01100100; | Outputs: P=%b | Expected: P=%d",
                 1967,
                 
                 P
                 , 
                 
                 20900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101011; B = 8'b00100100; // Expected: {'P': 6156}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101011; B = 8'b00100100; | Outputs: P=%b | Expected: P=%d",
                 1968,
                 
                 P
                 , 
                 
                 6156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011110; B = 8'b00000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011110; B = 8'b00000000; | Outputs: P=%b | Expected: P=%d",
                 1969,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001011; B = 8'b00000101; // Expected: {'P': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001011; B = 8'b00000101; | Outputs: P=%b | Expected: P=%d",
                 1970,
                 
                 P
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100000; B = 8'b11111101; // Expected: {'P': 8096}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100000; B = 8'b11111101; | Outputs: P=%b | Expected: P=%d",
                 1971,
                 
                 P
                 , 
                 
                 8096
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111000; B = 8'b00000011; // Expected: {'P': 168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111000; B = 8'b00000011; | Outputs: P=%b | Expected: P=%d",
                 1972,
                 
                 P
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110000; B = 8'b01000001; // Expected: {'P': 7280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110000; B = 8'b01000001; | Outputs: P=%b | Expected: P=%d",
                 1973,
                 
                 P
                 , 
                 
                 7280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010010; B = 8'b00001000; // Expected: {'P': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010010; B = 8'b00001000; | Outputs: P=%b | Expected: P=%d",
                 1974,
                 
                 P
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001001; B = 8'b00001001; // Expected: {'P': 81}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001001; B = 8'b00001001; | Outputs: P=%b | Expected: P=%d",
                 1975,
                 
                 P
                 , 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100010; B = 8'b00101010; // Expected: {'P': 4116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100010; B = 8'b00101010; | Outputs: P=%b | Expected: P=%d",
                 1976,
                 
                 P
                 , 
                 
                 4116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011100; B = 8'b11111001; // Expected: {'P': 6972}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011100; B = 8'b11111001; | Outputs: P=%b | Expected: P=%d",
                 1977,
                 
                 P
                 , 
                 
                 6972
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101001; B = 8'b10000000; // Expected: {'P': 21632}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101001; B = 8'b10000000; | Outputs: P=%b | Expected: P=%d",
                 1978,
                 
                 P
                 , 
                 
                 21632
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110100; B = 8'b01010001; // Expected: {'P': 19764}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110100; B = 8'b01010001; | Outputs: P=%b | Expected: P=%d",
                 1979,
                 
                 P
                 , 
                 
                 19764
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000011; B = 8'b01100000; // Expected: {'P': 12576}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000011; B = 8'b01100000; | Outputs: P=%b | Expected: P=%d",
                 1980,
                 
                 P
                 , 
                 
                 12576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100101; B = 8'b01001110; // Expected: {'P': 2886}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100101; B = 8'b01001110; | Outputs: P=%b | Expected: P=%d",
                 1981,
                 
                 P
                 , 
                 
                 2886
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110001; B = 8'b00101111; // Expected: {'P': 5311}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110001; B = 8'b00101111; | Outputs: P=%b | Expected: P=%d",
                 1982,
                 
                 P
                 , 
                 
                 5311
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100000; B = 8'b10111100; // Expected: {'P': 30080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100000; B = 8'b10111100; | Outputs: P=%b | Expected: P=%d",
                 1983,
                 
                 P
                 , 
                 
                 30080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111100; B = 8'b00110011; // Expected: {'P': 3060}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111100; B = 8'b00110011; | Outputs: P=%b | Expected: P=%d",
                 1984,
                 
                 P
                 , 
                 
                 3060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111110; B = 8'b01110100; // Expected: {'P': 22040}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111110; B = 8'b01110100; | Outputs: P=%b | Expected: P=%d",
                 1985,
                 
                 P
                 , 
                 
                 22040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010011; B = 8'b01000001; // Expected: {'P': 13715}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010011; B = 8'b01000001; | Outputs: P=%b | Expected: P=%d",
                 1986,
                 
                 P
                 , 
                 
                 13715
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000111; B = 8'b11110011; // Expected: {'P': 48357}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000111; B = 8'b11110011; | Outputs: P=%b | Expected: P=%d",
                 1987,
                 
                 P
                 , 
                 
                 48357
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101111; B = 8'b11101010; // Expected: {'P': 40950}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101111; B = 8'b11101010; | Outputs: P=%b | Expected: P=%d",
                 1988,
                 
                 P
                 , 
                 
                 40950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100100; B = 8'b10100110; // Expected: {'P': 37848}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100100; B = 8'b10100110; | Outputs: P=%b | Expected: P=%d",
                 1989,
                 
                 P
                 , 
                 
                 37848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110000; B = 8'b11100101; // Expected: {'P': 54960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110000; B = 8'b11100101; | Outputs: P=%b | Expected: P=%d",
                 1990,
                 
                 P
                 , 
                 
                 54960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001001; B = 8'b10110000; // Expected: {'P': 12848}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001001; B = 8'b10110000; | Outputs: P=%b | Expected: P=%d",
                 1991,
                 
                 P
                 , 
                 
                 12848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111011; B = 8'b11110111; // Expected: {'P': 14573}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111011; B = 8'b11110111; | Outputs: P=%b | Expected: P=%d",
                 1992,
                 
                 P
                 , 
                 
                 14573
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100111; B = 8'b10110100; // Expected: {'P': 7020}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100111; B = 8'b10110100; | Outputs: P=%b | Expected: P=%d",
                 1993,
                 
                 P
                 , 
                 
                 7020
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100110; B = 8'b10110110; // Expected: {'P': 30212}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100110; B = 8'b10110110; | Outputs: P=%b | Expected: P=%d",
                 1994,
                 
                 P
                 , 
                 
                 30212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111101; B = 8'b00011111; // Expected: {'P': 7843}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111101; B = 8'b00011111; | Outputs: P=%b | Expected: P=%d",
                 1995,
                 
                 P
                 , 
                 
                 7843
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010001; B = 8'b10000000; // Expected: {'P': 2176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010001; B = 8'b10000000; | Outputs: P=%b | Expected: P=%d",
                 1996,
                 
                 P
                 , 
                 
                 2176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110101; B = 8'b01111000; // Expected: {'P': 21720}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110101; B = 8'b01111000; | Outputs: P=%b | Expected: P=%d",
                 1997,
                 
                 P
                 , 
                 
                 21720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111000; B = 8'b11111000; // Expected: {'P': 61504}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111000; B = 8'b11111000; | Outputs: P=%b | Expected: P=%d",
                 1998,
                 
                 P
                 , 
                 
                 61504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011010; B = 8'b10000101; // Expected: {'P': 3458}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011010; B = 8'b10000101; | Outputs: P=%b | Expected: P=%d",
                 1999,
                 
                 P
                 , 
                 
                 3458
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100010; B = 8'b11001000; // Expected: {'P': 6800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100010; B = 8'b11001000; | Outputs: P=%b | Expected: P=%d",
                 2000,
                 
                 P
                 , 
                 
                 6800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101100; B = 8'b00001001; // Expected: {'P': 1548}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101100; B = 8'b00001001; | Outputs: P=%b | Expected: P=%d",
                 2001,
                 
                 P
                 , 
                 
                 1548
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101110; B = 8'b11000001; // Expected: {'P': 8878}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101110; B = 8'b11000001; | Outputs: P=%b | Expected: P=%d",
                 2002,
                 
                 P
                 , 
                 
                 8878
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100000; B = 8'b11011101; // Expected: {'P': 21216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100000; B = 8'b11011101; | Outputs: P=%b | Expected: P=%d",
                 2003,
                 
                 P
                 , 
                 
                 21216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110100; B = 8'b10110111; // Expected: {'P': 44652}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110100; B = 8'b10110111; | Outputs: P=%b | Expected: P=%d",
                 2004,
                 
                 P
                 , 
                 
                 44652
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011101; B = 8'b01010100; // Expected: {'P': 2436}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011101; B = 8'b01010100; | Outputs: P=%b | Expected: P=%d",
                 2005,
                 
                 P
                 , 
                 
                 2436
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010001; B = 8'b00000101; // Expected: {'P': 1045}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010001; B = 8'b00000101; | Outputs: P=%b | Expected: P=%d",
                 2006,
                 
                 P
                 , 
                 
                 1045
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001110; B = 8'b10100001; // Expected: {'P': 12558}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001110; B = 8'b10100001; | Outputs: P=%b | Expected: P=%d",
                 2007,
                 
                 P
                 , 
                 
                 12558
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010110; B = 8'b10000110; // Expected: {'P': 2948}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010110; B = 8'b10000110; | Outputs: P=%b | Expected: P=%d",
                 2008,
                 
                 P
                 , 
                 
                 2948
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001110; B = 8'b10000001; // Expected: {'P': 18318}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001110; B = 8'b10000001; | Outputs: P=%b | Expected: P=%d",
                 2009,
                 
                 P
                 , 
                 
                 18318
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011100; B = 8'b10000000; // Expected: {'P': 19968}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011100; B = 8'b10000000; | Outputs: P=%b | Expected: P=%d",
                 2010,
                 
                 P
                 , 
                 
                 19968
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111001; B = 8'b01101110; // Expected: {'P': 6270}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111001; B = 8'b01101110; | Outputs: P=%b | Expected: P=%d",
                 2011,
                 
                 P
                 , 
                 
                 6270
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100110; B = 8'b00110100; // Expected: {'P': 5304}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100110; B = 8'b00110100; | Outputs: P=%b | Expected: P=%d",
                 2012,
                 
                 P
                 , 
                 
                 5304
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000001; B = 8'b10110000; // Expected: {'P': 11440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000001; B = 8'b10110000; | Outputs: P=%b | Expected: P=%d",
                 2013,
                 
                 P
                 , 
                 
                 11440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101010; B = 8'b11101101; // Expected: {'P': 25122}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101010; B = 8'b11101101; | Outputs: P=%b | Expected: P=%d",
                 2014,
                 
                 P
                 , 
                 
                 25122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010001; B = 8'b10100011; // Expected: {'P': 2771}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010001; B = 8'b10100011; | Outputs: P=%b | Expected: P=%d",
                 2015,
                 
                 P
                 , 
                 
                 2771
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001000; B = 8'b11101010; // Expected: {'P': 31824}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001000; B = 8'b11101010; | Outputs: P=%b | Expected: P=%d",
                 2016,
                 
                 P
                 , 
                 
                 31824
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110000; B = 8'b00110110; // Expected: {'P': 12960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110000; B = 8'b00110110; | Outputs: P=%b | Expected: P=%d",
                 2017,
                 
                 P
                 , 
                 
                 12960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101011; B = 8'b01011101; // Expected: {'P': 15903}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101011; B = 8'b01011101; | Outputs: P=%b | Expected: P=%d",
                 2018,
                 
                 P
                 , 
                 
                 15903
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001101; B = 8'b10011101; // Expected: {'P': 32185}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001101; B = 8'b10011101; | Outputs: P=%b | Expected: P=%d",
                 2019,
                 
                 P
                 , 
                 
                 32185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000100; B = 8'b01101011; // Expected: {'P': 14124}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000100; B = 8'b01101011; | Outputs: P=%b | Expected: P=%d",
                 2020,
                 
                 P
                 , 
                 
                 14124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100101; B = 8'b00101110; // Expected: {'P': 10534}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100101; B = 8'b00101110; | Outputs: P=%b | Expected: P=%d",
                 2021,
                 
                 P
                 , 
                 
                 10534
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101100; B = 8'b11011011; // Expected: {'P': 51684}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101100; B = 8'b11011011; | Outputs: P=%b | Expected: P=%d",
                 2022,
                 
                 P
                 , 
                 
                 51684
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001000; B = 8'b10000011; // Expected: {'P': 17816}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001000; B = 8'b10000011; | Outputs: P=%b | Expected: P=%d",
                 2023,
                 
                 P
                 , 
                 
                 17816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101101; B = 8'b11101000; // Expected: {'P': 25288}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101101; B = 8'b11101000; | Outputs: P=%b | Expected: P=%d",
                 2024,
                 
                 P
                 , 
                 
                 25288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000100; B = 8'b00111010; // Expected: {'P': 11368}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000100; B = 8'b00111010; | Outputs: P=%b | Expected: P=%d",
                 2025,
                 
                 P
                 , 
                 
                 11368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100001; B = 8'b10100000; // Expected: {'P': 5280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100001; B = 8'b10100000; | Outputs: P=%b | Expected: P=%d",
                 2026,
                 
                 P
                 , 
                 
                 5280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111110; B = 8'b10011111; // Expected: {'P': 9858}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111110; B = 8'b10011111; | Outputs: P=%b | Expected: P=%d",
                 2027,
                 
                 P
                 , 
                 
                 9858
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111010; B = 8'b01101101; // Expected: {'P': 27250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111010; B = 8'b01101101; | Outputs: P=%b | Expected: P=%d",
                 2028,
                 
                 P
                 , 
                 
                 27250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010010; B = 8'b10100001; // Expected: {'P': 33810}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010010; B = 8'b10100001; | Outputs: P=%b | Expected: P=%d",
                 2029,
                 
                 P
                 , 
                 
                 33810
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111001; B = 8'b10111000; // Expected: {'P': 45816}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111001; B = 8'b10111000; | Outputs: P=%b | Expected: P=%d",
                 2030,
                 
                 P
                 , 
                 
                 45816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100110; B = 8'b11101000; // Expected: {'P': 8816}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100110; B = 8'b11101000; | Outputs: P=%b | Expected: P=%d",
                 2031,
                 
                 P
                 , 
                 
                 8816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110001; B = 8'b10011010; // Expected: {'P': 27258}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110001; B = 8'b10011010; | Outputs: P=%b | Expected: P=%d",
                 2032,
                 
                 P
                 , 
                 
                 27258
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101111; B = 8'b10101010; // Expected: {'P': 7990}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101111; B = 8'b10101010; | Outputs: P=%b | Expected: P=%d",
                 2033,
                 
                 P
                 , 
                 
                 7990
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011100; B = 8'b10100001; // Expected: {'P': 25116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011100; B = 8'b10100001; | Outputs: P=%b | Expected: P=%d",
                 2034,
                 
                 P
                 , 
                 
                 25116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011101; B = 8'b00011110; // Expected: {'P': 6630}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011101; B = 8'b00011110; | Outputs: P=%b | Expected: P=%d",
                 2035,
                 
                 P
                 , 
                 
                 6630
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100000; B = 8'b11100101; // Expected: {'P': 21984}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100000; B = 8'b11100101; | Outputs: P=%b | Expected: P=%d",
                 2036,
                 
                 P
                 , 
                 
                 21984
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011100; B = 8'b00000101; // Expected: {'P': 1100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011100; B = 8'b00000101; | Outputs: P=%b | Expected: P=%d",
                 2037,
                 
                 P
                 , 
                 
                 1100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101101; B = 8'b10011001; // Expected: {'P': 6885}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101101; B = 8'b10011001; | Outputs: P=%b | Expected: P=%d",
                 2038,
                 
                 P
                 , 
                 
                 6885
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000100; B = 8'b01000001; // Expected: {'P': 260}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000100; B = 8'b01000001; | Outputs: P=%b | Expected: P=%d",
                 2039,
                 
                 P
                 , 
                 
                 260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111101; B = 8'b10001001; // Expected: {'P': 34661}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111101; B = 8'b10001001; | Outputs: P=%b | Expected: P=%d",
                 2040,
                 
                 P
                 , 
                 
                 34661
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100101; B = 8'b00010011; // Expected: {'P': 3135}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100101; B = 8'b00010011; | Outputs: P=%b | Expected: P=%d",
                 2041,
                 
                 P
                 , 
                 
                 3135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110110; B = 8'b00110100; // Expected: {'P': 2808}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110110; B = 8'b00110100; | Outputs: P=%b | Expected: P=%d",
                 2042,
                 
                 P
                 , 
                 
                 2808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001000; B = 8'b00101011; // Expected: {'P': 5848}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001000; B = 8'b00101011; | Outputs: P=%b | Expected: P=%d",
                 2043,
                 
                 P
                 , 
                 
                 5848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001000; B = 8'b10000101; // Expected: {'P': 18088}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001000; B = 8'b10000101; | Outputs: P=%b | Expected: P=%d",
                 2044,
                 
                 P
                 , 
                 
                 18088
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011010; B = 8'b11001010; // Expected: {'P': 31108}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011010; B = 8'b11001010; | Outputs: P=%b | Expected: P=%d",
                 2045,
                 
                 P
                 , 
                 
                 31108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001100; B = 8'b10111110; // Expected: {'P': 26600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001100; B = 8'b10111110; | Outputs: P=%b | Expected: P=%d",
                 2046,
                 
                 P
                 , 
                 
                 26600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101010; B = 8'b00100100; // Expected: {'P': 3816}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101010; B = 8'b00100100; | Outputs: P=%b | Expected: P=%d",
                 2047,
                 
                 P
                 , 
                 
                 3816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111001; B = 8'b11000111; // Expected: {'P': 11343}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111001; B = 8'b11000111; | Outputs: P=%b | Expected: P=%d",
                 2048,
                 
                 P
                 , 
                 
                 11343
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001111; B = 8'b00000100; // Expected: {'P': 828}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001111; B = 8'b00000100; | Outputs: P=%b | Expected: P=%d",
                 2049,
                 
                 P
                 , 
                 
                 828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001110; B = 8'b10001010; // Expected: {'P': 10764}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001110; B = 8'b10001010; | Outputs: P=%b | Expected: P=%d",
                 2050,
                 
                 P
                 , 
                 
                 10764
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100110; B = 8'b01110010; // Expected: {'P': 4332}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100110; B = 8'b01110010; | Outputs: P=%b | Expected: P=%d",
                 2051,
                 
                 P
                 , 
                 
                 4332
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111010; B = 8'b11101100; // Expected: {'P': 43896}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111010; B = 8'b11101100; | Outputs: P=%b | Expected: P=%d",
                 2052,
                 
                 P
                 , 
                 
                 43896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000001; B = 8'b11001001; // Expected: {'P': 201}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000001; B = 8'b11001001; | Outputs: P=%b | Expected: P=%d",
                 2053,
                 
                 P
                 , 
                 
                 201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011010; B = 8'b11111001; // Expected: {'P': 38346}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011010; B = 8'b11111001; | Outputs: P=%b | Expected: P=%d",
                 2054,
                 
                 P
                 , 
                 
                 38346
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100000; B = 8'b10110110; // Expected: {'P': 29120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100000; B = 8'b10110110; | Outputs: P=%b | Expected: P=%d",
                 2055,
                 
                 P
                 , 
                 
                 29120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000000; B = 8'b01000100; // Expected: {'P': 8704}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000000; B = 8'b01000100; | Outputs: P=%b | Expected: P=%d",
                 2056,
                 
                 P
                 , 
                 
                 8704
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001000; B = 8'b10110111; // Expected: {'P': 1464}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001000; B = 8'b10110111; | Outputs: P=%b | Expected: P=%d",
                 2057,
                 
                 P
                 , 
                 
                 1464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010110; B = 8'b10100001; // Expected: {'P': 3542}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010110; B = 8'b10100001; | Outputs: P=%b | Expected: P=%d",
                 2058,
                 
                 P
                 , 
                 
                 3542
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110110; B = 8'b10101000; // Expected: {'P': 41328}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110110; B = 8'b10101000; | Outputs: P=%b | Expected: P=%d",
                 2059,
                 
                 P
                 , 
                 
                 41328
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101100; B = 8'b10010011; // Expected: {'P': 15876}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101100; B = 8'b10010011; | Outputs: P=%b | Expected: P=%d",
                 2060,
                 
                 P
                 , 
                 
                 15876
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011111; B = 8'b11010000; // Expected: {'P': 6448}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011111; B = 8'b11010000; | Outputs: P=%b | Expected: P=%d",
                 2061,
                 
                 P
                 , 
                 
                 6448
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111000; B = 8'b01010101; // Expected: {'P': 15640}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111000; B = 8'b01010101; | Outputs: P=%b | Expected: P=%d",
                 2062,
                 
                 P
                 , 
                 
                 15640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100010; B = 8'b01010010; // Expected: {'P': 8036}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100010; B = 8'b01010010; | Outputs: P=%b | Expected: P=%d",
                 2063,
                 
                 P
                 , 
                 
                 8036
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101101; B = 8'b01111010; // Expected: {'P': 28914}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101101; B = 8'b01111010; | Outputs: P=%b | Expected: P=%d",
                 2064,
                 
                 P
                 , 
                 
                 28914
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110110; B = 8'b10100000; // Expected: {'P': 29120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110110; B = 8'b10100000; | Outputs: P=%b | Expected: P=%d",
                 2065,
                 
                 P
                 , 
                 
                 29120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111000; B = 8'b00111010; // Expected: {'P': 3248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111000; B = 8'b00111010; | Outputs: P=%b | Expected: P=%d",
                 2066,
                 
                 P
                 , 
                 
                 3248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011000; B = 8'b01110010; // Expected: {'P': 2736}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011000; B = 8'b01110010; | Outputs: P=%b | Expected: P=%d",
                 2067,
                 
                 P
                 , 
                 
                 2736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010010; B = 8'b00110000; // Expected: {'P': 7008}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010010; B = 8'b00110000; | Outputs: P=%b | Expected: P=%d",
                 2068,
                 
                 P
                 , 
                 
                 7008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000001; B = 8'b10011000; // Expected: {'P': 19608}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000001; B = 8'b10011000; | Outputs: P=%b | Expected: P=%d",
                 2069,
                 
                 P
                 , 
                 
                 19608
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101100; B = 8'b11110101; // Expected: {'P': 42140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101100; B = 8'b11110101; | Outputs: P=%b | Expected: P=%d",
                 2070,
                 
                 P
                 , 
                 
                 42140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111111; B = 8'b11000101; // Expected: {'P': 12411}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111111; B = 8'b11000101; | Outputs: P=%b | Expected: P=%d",
                 2071,
                 
                 P
                 , 
                 
                 12411
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100100; B = 8'b00111000; // Expected: {'P': 9184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100100; B = 8'b00111000; | Outputs: P=%b | Expected: P=%d",
                 2072,
                 
                 P
                 , 
                 
                 9184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101011; B = 8'b11000010; // Expected: {'P': 33174}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101011; B = 8'b11000010; | Outputs: P=%b | Expected: P=%d",
                 2073,
                 
                 P
                 , 
                 
                 33174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010001; B = 8'b00110011; // Expected: {'P': 4131}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010001; B = 8'b00110011; | Outputs: P=%b | Expected: P=%d",
                 2074,
                 
                 P
                 , 
                 
                 4131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101010; B = 8'b00101100; // Expected: {'P': 4664}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101010; B = 8'b00101100; | Outputs: P=%b | Expected: P=%d",
                 2075,
                 
                 P
                 , 
                 
                 4664
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110010; B = 8'b01100000; // Expected: {'P': 4800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110010; B = 8'b01100000; | Outputs: P=%b | Expected: P=%d",
                 2076,
                 
                 P
                 , 
                 
                 4800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010000; B = 8'b01110101; // Expected: {'P': 1872}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010000; B = 8'b01110101; | Outputs: P=%b | Expected: P=%d",
                 2077,
                 
                 P
                 , 
                 
                 1872
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001100; B = 8'b00010001; // Expected: {'P': 2380}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001100; B = 8'b00010001; | Outputs: P=%b | Expected: P=%d",
                 2078,
                 
                 P
                 , 
                 
                 2380
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011101; B = 8'b00000010; // Expected: {'P': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011101; B = 8'b00000010; | Outputs: P=%b | Expected: P=%d",
                 2079,
                 
                 P
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000000; B = 8'b00101001; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000000; B = 8'b00101001; | Outputs: P=%b | Expected: P=%d",
                 2080,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101101; B = 8'b00000010; // Expected: {'P': 474}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101101; B = 8'b00000010; | Outputs: P=%b | Expected: P=%d",
                 2081,
                 
                 P
                 , 
                 
                 474
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100110; B = 8'b00101110; // Expected: {'P': 7636}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100110; B = 8'b00101110; | Outputs: P=%b | Expected: P=%d",
                 2082,
                 
                 P
                 , 
                 
                 7636
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101011; B = 8'b00001110; // Expected: {'P': 1498}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101011; B = 8'b00001110; | Outputs: P=%b | Expected: P=%d",
                 2083,
                 
                 P
                 , 
                 
                 1498
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101001; B = 8'b01100001; // Expected: {'P': 22601}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101001; B = 8'b01100001; | Outputs: P=%b | Expected: P=%d",
                 2084,
                 
                 P
                 , 
                 
                 22601
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101110; B = 8'b01000010; // Expected: {'P': 15708}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101110; B = 8'b01000010; | Outputs: P=%b | Expected: P=%d",
                 2085,
                 
                 P
                 , 
                 
                 15708
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101110; B = 8'b01010001; // Expected: {'P': 19278}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101110; B = 8'b01010001; | Outputs: P=%b | Expected: P=%d",
                 2086,
                 
                 P
                 , 
                 
                 19278
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101101; B = 8'b11001101; // Expected: {'P': 22345}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101101; B = 8'b11001101; | Outputs: P=%b | Expected: P=%d",
                 2087,
                 
                 P
                 , 
                 
                 22345
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010101; B = 8'b01111111; // Expected: {'P': 10795}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010101; B = 8'b01111111; | Outputs: P=%b | Expected: P=%d",
                 2088,
                 
                 P
                 , 
                 
                 10795
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101011; B = 8'b10001111; // Expected: {'P': 15301}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101011; B = 8'b10001111; | Outputs: P=%b | Expected: P=%d",
                 2089,
                 
                 P
                 , 
                 
                 15301
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110101; B = 8'b01111100; // Expected: {'P': 22444}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110101; B = 8'b01111100; | Outputs: P=%b | Expected: P=%d",
                 2090,
                 
                 P
                 , 
                 
                 22444
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101110; B = 8'b11101101; // Expected: {'P': 26070}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101110; B = 8'b11101101; | Outputs: P=%b | Expected: P=%d",
                 2091,
                 
                 P
                 , 
                 
                 26070
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011000; B = 8'b00010000; // Expected: {'P': 3456}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011000; B = 8'b00010000; | Outputs: P=%b | Expected: P=%d",
                 2092,
                 
                 P
                 , 
                 
                 3456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011010; B = 8'b10100110; // Expected: {'P': 14940}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011010; B = 8'b10100110; | Outputs: P=%b | Expected: P=%d",
                 2093,
                 
                 P
                 , 
                 
                 14940
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100100; B = 8'b01011111; // Expected: {'P': 15580}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100100; B = 8'b01011111; | Outputs: P=%b | Expected: P=%d",
                 2094,
                 
                 P
                 , 
                 
                 15580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001111; B = 8'b00110000; // Expected: {'P': 6864}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001111; B = 8'b00110000; | Outputs: P=%b | Expected: P=%d",
                 2095,
                 
                 P
                 , 
                 
                 6864
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100011; B = 8'b00111001; // Expected: {'P': 1995}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100011; B = 8'b00111001; | Outputs: P=%b | Expected: P=%d",
                 2096,
                 
                 P
                 , 
                 
                 1995
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011100; B = 8'b00100010; // Expected: {'P': 952}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011100; B = 8'b00100010; | Outputs: P=%b | Expected: P=%d",
                 2097,
                 
                 P
                 , 
                 
                 952
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001001; B = 8'b01110101; // Expected: {'P': 23517}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001001; B = 8'b01110101; | Outputs: P=%b | Expected: P=%d",
                 2098,
                 
                 P
                 , 
                 
                 23517
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000000; B = 8'b11110110; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000000; B = 8'b11110110; | Outputs: P=%b | Expected: P=%d",
                 2099,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001011; B = 8'b00111011; // Expected: {'P': 11977}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001011; B = 8'b00111011; | Outputs: P=%b | Expected: P=%d",
                 2100,
                 
                 P
                 , 
                 
                 11977
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100010; B = 8'b00100001; // Expected: {'P': 5346}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100010; B = 8'b00100001; | Outputs: P=%b | Expected: P=%d",
                 2101,
                 
                 P
                 , 
                 
                 5346
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111001; B = 8'b11011011; // Expected: {'P': 54531}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111001; B = 8'b11011011; | Outputs: P=%b | Expected: P=%d",
                 2102,
                 
                 P
                 , 
                 
                 54531
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001011; B = 8'b10101001; // Expected: {'P': 23491}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001011; B = 8'b10101001; | Outputs: P=%b | Expected: P=%d",
                 2103,
                 
                 P
                 , 
                 
                 23491
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001000; B = 8'b00100101; // Expected: {'P': 296}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001000; B = 8'b00100101; | Outputs: P=%b | Expected: P=%d",
                 2104,
                 
                 P
                 , 
                 
                 296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110000; B = 8'b00100110; // Expected: {'P': 6688}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110000; B = 8'b00100110; | Outputs: P=%b | Expected: P=%d",
                 2105,
                 
                 P
                 , 
                 
                 6688
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011011; B = 8'b10011010; // Expected: {'P': 23870}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011011; B = 8'b10011010; | Outputs: P=%b | Expected: P=%d",
                 2106,
                 
                 P
                 , 
                 
                 23870
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100100; B = 8'b10001001; // Expected: {'P': 13700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100100; B = 8'b10001001; | Outputs: P=%b | Expected: P=%d",
                 2107,
                 
                 P
                 , 
                 
                 13700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011010; B = 8'b11100010; // Expected: {'P': 34804}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011010; B = 8'b11100010; | Outputs: P=%b | Expected: P=%d",
                 2108,
                 
                 P
                 , 
                 
                 34804
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100000; B = 8'b00011110; // Expected: {'P': 6720}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100000; B = 8'b00011110; | Outputs: P=%b | Expected: P=%d",
                 2109,
                 
                 P
                 , 
                 
                 6720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000100; B = 8'b01000100; // Expected: {'P': 13328}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000100; B = 8'b01000100; | Outputs: P=%b | Expected: P=%d",
                 2110,
                 
                 P
                 , 
                 
                 13328
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100101; B = 8'b01100000; // Expected: {'P': 3552}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100101; B = 8'b01100000; | Outputs: P=%b | Expected: P=%d",
                 2111,
                 
                 P
                 , 
                 
                 3552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000010; B = 8'b01000011; // Expected: {'P': 8710}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000010; B = 8'b01000011; | Outputs: P=%b | Expected: P=%d",
                 2112,
                 
                 P
                 , 
                 
                 8710
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101110; B = 8'b10100100; // Expected: {'P': 18040}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101110; B = 8'b10100100; | Outputs: P=%b | Expected: P=%d",
                 2113,
                 
                 P
                 , 
                 
                 18040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010100; B = 8'b01001110; // Expected: {'P': 11544}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010100; B = 8'b01001110; | Outputs: P=%b | Expected: P=%d",
                 2114,
                 
                 P
                 , 
                 
                 11544
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100001; B = 8'b01010001; // Expected: {'P': 7857}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100001; B = 8'b01010001; | Outputs: P=%b | Expected: P=%d",
                 2115,
                 
                 P
                 , 
                 
                 7857
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100010; B = 8'b00010111; // Expected: {'P': 5198}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100010; B = 8'b00010111; | Outputs: P=%b | Expected: P=%d",
                 2116,
                 
                 P
                 , 
                 
                 5198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010001; B = 8'b11110101; // Expected: {'P': 51205}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010001; B = 8'b11110101; | Outputs: P=%b | Expected: P=%d",
                 2117,
                 
                 P
                 , 
                 
                 51205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100010; B = 8'b01001010; // Expected: {'P': 7252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100010; B = 8'b01001010; | Outputs: P=%b | Expected: P=%d",
                 2118,
                 
                 P
                 , 
                 
                 7252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010110; B = 8'b00010101; // Expected: {'P': 462}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010110; B = 8'b00010101; | Outputs: P=%b | Expected: P=%d",
                 2119,
                 
                 P
                 , 
                 
                 462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001101; B = 8'b10110100; // Expected: {'P': 25380}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001101; B = 8'b10110100; | Outputs: P=%b | Expected: P=%d",
                 2120,
                 
                 P
                 , 
                 
                 25380
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101011; B = 8'b10001001; // Expected: {'P': 32195}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101011; B = 8'b10001001; | Outputs: P=%b | Expected: P=%d",
                 2121,
                 
                 P
                 , 
                 
                 32195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011000; B = 8'b00110010; // Expected: {'P': 1200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011000; B = 8'b00110010; | Outputs: P=%b | Expected: P=%d",
                 2122,
                 
                 P
                 , 
                 
                 1200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011010; B = 8'b00111001; // Expected: {'P': 12426}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011010; B = 8'b00111001; | Outputs: P=%b | Expected: P=%d",
                 2123,
                 
                 P
                 , 
                 
                 12426
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100100; B = 8'b00010111; // Expected: {'P': 2300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100100; B = 8'b00010111; | Outputs: P=%b | Expected: P=%d",
                 2124,
                 
                 P
                 , 
                 
                 2300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001011; B = 8'b10101100; // Expected: {'P': 23908}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001011; B = 8'b10101100; | Outputs: P=%b | Expected: P=%d",
                 2125,
                 
                 P
                 , 
                 
                 23908
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110011; B = 8'b00111111; // Expected: {'P': 15309}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110011; B = 8'b00111111; | Outputs: P=%b | Expected: P=%d",
                 2126,
                 
                 P
                 , 
                 
                 15309
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111011; B = 8'b10100010; // Expected: {'P': 9558}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111011; B = 8'b10100010; | Outputs: P=%b | Expected: P=%d",
                 2127,
                 
                 P
                 , 
                 
                 9558
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001100; B = 8'b11011010; // Expected: {'P': 44472}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001100; B = 8'b11011010; | Outputs: P=%b | Expected: P=%d",
                 2128,
                 
                 P
                 , 
                 
                 44472
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000100; B = 8'b00000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000100; B = 8'b00000000; | Outputs: P=%b | Expected: P=%d",
                 2129,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111001; B = 8'b01000001; // Expected: {'P': 16185}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111001; B = 8'b01000001; | Outputs: P=%b | Expected: P=%d",
                 2130,
                 
                 P
                 , 
                 
                 16185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000100; B = 8'b00001110; // Expected: {'P': 1848}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000100; B = 8'b00001110; | Outputs: P=%b | Expected: P=%d",
                 2131,
                 
                 P
                 , 
                 
                 1848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110011; B = 8'b00100011; // Expected: {'P': 4025}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110011; B = 8'b00100011; | Outputs: P=%b | Expected: P=%d",
                 2132,
                 
                 P
                 , 
                 
                 4025
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001000; B = 8'b10111100; // Expected: {'P': 1504}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001000; B = 8'b10111100; | Outputs: P=%b | Expected: P=%d",
                 2133,
                 
                 P
                 , 
                 
                 1504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100011; B = 8'b11100100; // Expected: {'P': 37164}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100011; B = 8'b11100100; | Outputs: P=%b | Expected: P=%d",
                 2134,
                 
                 P
                 , 
                 
                 37164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101011; B = 8'b00101110; // Expected: {'P': 1978}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101011; B = 8'b00101110; | Outputs: P=%b | Expected: P=%d",
                 2135,
                 
                 P
                 , 
                 
                 1978
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010011; B = 8'b01010000; // Expected: {'P': 16880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010011; B = 8'b01010000; | Outputs: P=%b | Expected: P=%d",
                 2136,
                 
                 P
                 , 
                 
                 16880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100010; B = 8'b00100010; // Expected: {'P': 1156}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100010; B = 8'b00100010; | Outputs: P=%b | Expected: P=%d",
                 2137,
                 
                 P
                 , 
                 
                 1156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000011; B = 8'b01100110; // Expected: {'P': 19890}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000011; B = 8'b01100110; | Outputs: P=%b | Expected: P=%d",
                 2138,
                 
                 P
                 , 
                 
                 19890
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000000; B = 8'b00100101; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000000; B = 8'b00100101; | Outputs: P=%b | Expected: P=%d",
                 2139,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011011; B = 8'b10011111; // Expected: {'P': 34821}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011011; B = 8'b10011111; | Outputs: P=%b | Expected: P=%d",
                 2140,
                 
                 P
                 , 
                 
                 34821
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100100; B = 8'b10011001; // Expected: {'P': 15300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100100; B = 8'b10011001; | Outputs: P=%b | Expected: P=%d",
                 2141,
                 
                 P
                 , 
                 
                 15300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110101; B = 8'b11101001; // Expected: {'P': 27261}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110101; B = 8'b11101001; | Outputs: P=%b | Expected: P=%d",
                 2142,
                 
                 P
                 , 
                 
                 27261
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111101; B = 8'b00000100; // Expected: {'P': 500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111101; B = 8'b00000100; | Outputs: P=%b | Expected: P=%d",
                 2143,
                 
                 P
                 , 
                 
                 500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110111; B = 8'b01111111; // Expected: {'P': 6985}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110111; B = 8'b01111111; | Outputs: P=%b | Expected: P=%d",
                 2144,
                 
                 P
                 , 
                 
                 6985
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010001; B = 8'b11010111; // Expected: {'P': 17415}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010001; B = 8'b11010111; | Outputs: P=%b | Expected: P=%d",
                 2145,
                 
                 P
                 , 
                 
                 17415
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001000; B = 8'b01100001; // Expected: {'P': 776}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001000; B = 8'b01100001; | Outputs: P=%b | Expected: P=%d",
                 2146,
                 
                 P
                 , 
                 
                 776
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001011; B = 8'b10010011; // Expected: {'P': 11025}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001011; B = 8'b10010011; | Outputs: P=%b | Expected: P=%d",
                 2147,
                 
                 P
                 , 
                 
                 11025
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010011; B = 8'b01000001; // Expected: {'P': 5395}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010011; B = 8'b01000001; | Outputs: P=%b | Expected: P=%d",
                 2148,
                 
                 P
                 , 
                 
                 5395
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110011; B = 8'b11011110; // Expected: {'P': 11322}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110011; B = 8'b11011110; | Outputs: P=%b | Expected: P=%d",
                 2149,
                 
                 P
                 , 
                 
                 11322
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001111; B = 8'b01010110; // Expected: {'P': 1290}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001111; B = 8'b01010110; | Outputs: P=%b | Expected: P=%d",
                 2150,
                 
                 P
                 , 
                 
                 1290
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001101; B = 8'b01011000; // Expected: {'P': 12408}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001101; B = 8'b01011000; | Outputs: P=%b | Expected: P=%d",
                 2151,
                 
                 P
                 , 
                 
                 12408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000000; B = 8'b10110011; // Expected: {'P': 22912}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000000; B = 8'b10110011; | Outputs: P=%b | Expected: P=%d",
                 2152,
                 
                 P
                 , 
                 
                 22912
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110001; B = 8'b01100011; // Expected: {'P': 17523}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110001; B = 8'b01100011; | Outputs: P=%b | Expected: P=%d",
                 2153,
                 
                 P
                 , 
                 
                 17523
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100010; B = 8'b00101111; // Expected: {'P': 1598}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100010; B = 8'b00101111; | Outputs: P=%b | Expected: P=%d",
                 2154,
                 
                 P
                 , 
                 
                 1598
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111101; B = 8'b10011111; // Expected: {'P': 19875}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111101; B = 8'b10011111; | Outputs: P=%b | Expected: P=%d",
                 2155,
                 
                 P
                 , 
                 
                 19875
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100100; B = 8'b01111011; // Expected: {'P': 4428}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100100; B = 8'b01111011; | Outputs: P=%b | Expected: P=%d",
                 2156,
                 
                 P
                 , 
                 
                 4428
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111101; B = 8'b01111111; // Expected: {'P': 7747}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111101; B = 8'b01111111; | Outputs: P=%b | Expected: P=%d",
                 2157,
                 
                 P
                 , 
                 
                 7747
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111011; B = 8'b11000101; // Expected: {'P': 11623}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111011; B = 8'b11000101; | Outputs: P=%b | Expected: P=%d",
                 2158,
                 
                 P
                 , 
                 
                 11623
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111110; B = 8'b00001000; // Expected: {'P': 1008}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111110; B = 8'b00001000; | Outputs: P=%b | Expected: P=%d",
                 2159,
                 
                 P
                 , 
                 
                 1008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010101; B = 8'b11001110; // Expected: {'P': 30694}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010101; B = 8'b11001110; | Outputs: P=%b | Expected: P=%d",
                 2160,
                 
                 P
                 , 
                 
                 30694
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110110; B = 8'b10011110; // Expected: {'P': 28756}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110110; B = 8'b10011110; | Outputs: P=%b | Expected: P=%d",
                 2161,
                 
                 P
                 , 
                 
                 28756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010101; B = 8'b10101011; // Expected: {'P': 25479}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010101; B = 8'b10101011; | Outputs: P=%b | Expected: P=%d",
                 2162,
                 
                 P
                 , 
                 
                 25479
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111000; B = 8'b00110111; // Expected: {'P': 10120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111000; B = 8'b00110111; | Outputs: P=%b | Expected: P=%d",
                 2163,
                 
                 P
                 , 
                 
                 10120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010100; B = 8'b01100000; // Expected: {'P': 1920}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010100; B = 8'b01100000; | Outputs: P=%b | Expected: P=%d",
                 2164,
                 
                 P
                 , 
                 
                 1920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110100; B = 8'b10010001; // Expected: {'P': 16820}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110100; B = 8'b10010001; | Outputs: P=%b | Expected: P=%d",
                 2165,
                 
                 P
                 , 
                 
                 16820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110011; B = 8'b01101001; // Expected: {'P': 18795}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110011; B = 8'b01101001; | Outputs: P=%b | Expected: P=%d",
                 2166,
                 
                 P
                 , 
                 
                 18795
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011110; B = 8'b11100110; // Expected: {'P': 51060}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011110; B = 8'b11100110; | Outputs: P=%b | Expected: P=%d",
                 2167,
                 
                 P
                 , 
                 
                 51060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001110; B = 8'b00111101; // Expected: {'P': 8662}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001110; B = 8'b00111101; | Outputs: P=%b | Expected: P=%d",
                 2168,
                 
                 P
                 , 
                 
                 8662
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011000; B = 8'b01010001; // Expected: {'P': 1944}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011000; B = 8'b01010001; | Outputs: P=%b | Expected: P=%d",
                 2169,
                 
                 P
                 , 
                 
                 1944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000001; B = 8'b11101000; // Expected: {'P': 15080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000001; B = 8'b11101000; | Outputs: P=%b | Expected: P=%d",
                 2170,
                 
                 P
                 , 
                 
                 15080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000000; B = 8'b00001100; // Expected: {'P': 2304}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000000; B = 8'b00001100; | Outputs: P=%b | Expected: P=%d",
                 2171,
                 
                 P
                 , 
                 
                 2304
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001001; B = 8'b00011111; // Expected: {'P': 6231}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001001; B = 8'b00011111; | Outputs: P=%b | Expected: P=%d",
                 2172,
                 
                 P
                 , 
                 
                 6231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111000; B = 8'b11110001; // Expected: {'P': 13496}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111000; B = 8'b11110001; | Outputs: P=%b | Expected: P=%d",
                 2173,
                 
                 P
                 , 
                 
                 13496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110001; B = 8'b00000011; // Expected: {'P': 147}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110001; B = 8'b00000011; | Outputs: P=%b | Expected: P=%d",
                 2174,
                 
                 P
                 , 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100011; B = 8'b11001011; // Expected: {'P': 7105}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100011; B = 8'b11001011; | Outputs: P=%b | Expected: P=%d",
                 2175,
                 
                 P
                 , 
                 
                 7105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111101; B = 8'b10111110; // Expected: {'P': 11590}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111101; B = 8'b10111110; | Outputs: P=%b | Expected: P=%d",
                 2176,
                 
                 P
                 , 
                 
                 11590
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101010; B = 8'b01111101; // Expected: {'P': 13250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101010; B = 8'b01111101; | Outputs: P=%b | Expected: P=%d",
                 2177,
                 
                 P
                 , 
                 
                 13250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001101; B = 8'b10011110; // Expected: {'P': 22278}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001101; B = 8'b10011110; | Outputs: P=%b | Expected: P=%d",
                 2178,
                 
                 P
                 , 
                 
                 22278
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001111; B = 8'b11000101; // Expected: {'P': 28171}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001111; B = 8'b11000101; | Outputs: P=%b | Expected: P=%d",
                 2179,
                 
                 P
                 , 
                 
                 28171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000011; B = 8'b01100101; // Expected: {'P': 6767}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000011; B = 8'b01100101; | Outputs: P=%b | Expected: P=%d",
                 2180,
                 
                 P
                 , 
                 
                 6767
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110001; B = 8'b01010001; // Expected: {'P': 14337}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110001; B = 8'b01010001; | Outputs: P=%b | Expected: P=%d",
                 2181,
                 
                 P
                 , 
                 
                 14337
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110101; B = 8'b01010101; // Expected: {'P': 9945}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110101; B = 8'b01010101; | Outputs: P=%b | Expected: P=%d",
                 2182,
                 
                 P
                 , 
                 
                 9945
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001010; B = 8'b00111110; // Expected: {'P': 8556}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001010; B = 8'b00111110; | Outputs: P=%b | Expected: P=%d",
                 2183,
                 
                 P
                 , 
                 
                 8556
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101100; B = 8'b01111010; // Expected: {'P': 5368}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101100; B = 8'b01111010; | Outputs: P=%b | Expected: P=%d",
                 2184,
                 
                 P
                 , 
                 
                 5368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001000; B = 8'b01001110; // Expected: {'P': 15600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001000; B = 8'b01001110; | Outputs: P=%b | Expected: P=%d",
                 2185,
                 
                 P
                 , 
                 
                 15600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110100; B = 8'b00000011; // Expected: {'P': 540}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110100; B = 8'b00000011; | Outputs: P=%b | Expected: P=%d",
                 2186,
                 
                 P
                 , 
                 
                 540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000001; B = 8'b00111000; // Expected: {'P': 10808}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000001; B = 8'b00111000; | Outputs: P=%b | Expected: P=%d",
                 2187,
                 
                 P
                 , 
                 
                 10808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010100; B = 8'b10111100; // Expected: {'P': 3760}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010100; B = 8'b10111100; | Outputs: P=%b | Expected: P=%d",
                 2188,
                 
                 P
                 , 
                 
                 3760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010110; B = 8'b11100110; // Expected: {'P': 34500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010110; B = 8'b11100110; | Outputs: P=%b | Expected: P=%d",
                 2189,
                 
                 P
                 , 
                 
                 34500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100111; B = 8'b10100110; // Expected: {'P': 17098}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100111; B = 8'b10100110; | Outputs: P=%b | Expected: P=%d",
                 2190,
                 
                 P
                 , 
                 
                 17098
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001111; B = 8'b01000111; // Expected: {'P': 1065}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001111; B = 8'b01000111; | Outputs: P=%b | Expected: P=%d",
                 2191,
                 
                 P
                 , 
                 
                 1065
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111110; B = 8'b01010010; // Expected: {'P': 15580}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111110; B = 8'b01010010; | Outputs: P=%b | Expected: P=%d",
                 2192,
                 
                 P
                 , 
                 
                 15580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110110; B = 8'b00010011; // Expected: {'P': 1026}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110110; B = 8'b00010011; | Outputs: P=%b | Expected: P=%d",
                 2193,
                 
                 P
                 , 
                 
                 1026
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010001; B = 8'b11000000; // Expected: {'P': 15552}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010001; B = 8'b11000000; | Outputs: P=%b | Expected: P=%d",
                 2194,
                 
                 P
                 , 
                 
                 15552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111001; B = 8'b01010100; // Expected: {'P': 15540}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111001; B = 8'b01010100; | Outputs: P=%b | Expected: P=%d",
                 2195,
                 
                 P
                 , 
                 
                 15540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001010; B = 8'b00110111; // Expected: {'P': 4070}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001010; B = 8'b00110111; | Outputs: P=%b | Expected: P=%d",
                 2196,
                 
                 P
                 , 
                 
                 4070
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011110; B = 8'b11000000; // Expected: {'P': 18048}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011110; B = 8'b11000000; | Outputs: P=%b | Expected: P=%d",
                 2197,
                 
                 P
                 , 
                 
                 18048
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101110; B = 8'b01010011; // Expected: {'P': 19754}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101110; B = 8'b01010011; | Outputs: P=%b | Expected: P=%d",
                 2198,
                 
                 P
                 , 
                 
                 19754
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000101; B = 8'b10001000; // Expected: {'P': 26792}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000101; B = 8'b10001000; | Outputs: P=%b | Expected: P=%d",
                 2199,
                 
                 P
                 , 
                 
                 26792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111100; B = 8'b01010010; // Expected: {'P': 4920}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111100; B = 8'b01010010; | Outputs: P=%b | Expected: P=%d",
                 2200,
                 
                 P
                 , 
                 
                 4920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110001; B = 8'b11011001; // Expected: {'P': 52297}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110001; B = 8'b11011001; | Outputs: P=%b | Expected: P=%d",
                 2201,
                 
                 P
                 , 
                 
                 52297
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000011; B = 8'b10000010; // Expected: {'P': 25350}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000011; B = 8'b10000010; | Outputs: P=%b | Expected: P=%d",
                 2202,
                 
                 P
                 , 
                 
                 25350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011000; B = 8'b01110100; // Expected: {'P': 2784}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011000; B = 8'b01110100; | Outputs: P=%b | Expected: P=%d",
                 2203,
                 
                 P
                 , 
                 
                 2784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101110; B = 8'b10011010; // Expected: {'P': 16940}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101110; B = 8'b10011010; | Outputs: P=%b | Expected: P=%d",
                 2204,
                 
                 P
                 , 
                 
                 16940
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100011; B = 8'b11110111; // Expected: {'P': 24453}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100011; B = 8'b11110111; | Outputs: P=%b | Expected: P=%d",
                 2205,
                 
                 P
                 , 
                 
                 24453
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101011; B = 8'b01111001; // Expected: {'P': 12947}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101011; B = 8'b01111001; | Outputs: P=%b | Expected: P=%d",
                 2206,
                 
                 P
                 , 
                 
                 12947
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010001; B = 8'b11010111; // Expected: {'P': 44935}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010001; B = 8'b11010111; | Outputs: P=%b | Expected: P=%d",
                 2207,
                 
                 P
                 , 
                 
                 44935
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010110; B = 8'b00000011; // Expected: {'P': 642}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010110; B = 8'b00000011; | Outputs: P=%b | Expected: P=%d",
                 2208,
                 
                 P
                 , 
                 
                 642
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101010; B = 8'b11010110; // Expected: {'P': 36380}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101010; B = 8'b11010110; | Outputs: P=%b | Expected: P=%d",
                 2209,
                 
                 P
                 , 
                 
                 36380
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110011; B = 8'b10110110; // Expected: {'P': 32578}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110011; B = 8'b10110110; | Outputs: P=%b | Expected: P=%d",
                 2210,
                 
                 P
                 , 
                 
                 32578
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010001; B = 8'b00011111; // Expected: {'P': 6479}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010001; B = 8'b00011111; | Outputs: P=%b | Expected: P=%d",
                 2211,
                 
                 P
                 , 
                 
                 6479
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000010; B = 8'b11011000; // Expected: {'P': 432}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000010; B = 8'b11011000; | Outputs: P=%b | Expected: P=%d",
                 2212,
                 
                 P
                 , 
                 
                 432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110000; B = 8'b01110101; // Expected: {'P': 20592}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110000; B = 8'b01110101; | Outputs: P=%b | Expected: P=%d",
                 2213,
                 
                 P
                 , 
                 
                 20592
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010000; B = 8'b11010010; // Expected: {'P': 16800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010000; B = 8'b11010010; | Outputs: P=%b | Expected: P=%d",
                 2214,
                 
                 P
                 , 
                 
                 16800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001011; B = 8'b01010101; // Expected: {'P': 6375}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001011; B = 8'b01010101; | Outputs: P=%b | Expected: P=%d",
                 2215,
                 
                 P
                 , 
                 
                 6375
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001000; B = 8'b11001000; // Expected: {'P': 27200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001000; B = 8'b11001000; | Outputs: P=%b | Expected: P=%d",
                 2216,
                 
                 P
                 , 
                 
                 27200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001001; B = 8'b10010101; // Expected: {'P': 1341}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001001; B = 8'b10010101; | Outputs: P=%b | Expected: P=%d",
                 2217,
                 
                 P
                 , 
                 
                 1341
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100111; B = 8'b10010011; // Expected: {'P': 15141}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100111; B = 8'b10010011; | Outputs: P=%b | Expected: P=%d",
                 2218,
                 
                 P
                 , 
                 
                 15141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100101; B = 8'b00001100; // Expected: {'P': 1980}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100101; B = 8'b00001100; | Outputs: P=%b | Expected: P=%d",
                 2219,
                 
                 P
                 , 
                 
                 1980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001001; B = 8'b11011000; // Expected: {'P': 1944}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001001; B = 8'b11011000; | Outputs: P=%b | Expected: P=%d",
                 2220,
                 
                 P
                 , 
                 
                 1944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000101; B = 8'b00110011; // Expected: {'P': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000101; B = 8'b00110011; | Outputs: P=%b | Expected: P=%d",
                 2221,
                 
                 P
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100011; B = 8'b00101000; // Expected: {'P': 1400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100011; B = 8'b00101000; | Outputs: P=%b | Expected: P=%d",
                 2222,
                 
                 P
                 , 
                 
                 1400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010101; B = 8'b00001101; // Expected: {'P': 273}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010101; B = 8'b00001101; | Outputs: P=%b | Expected: P=%d",
                 2223,
                 
                 P
                 , 
                 
                 273
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010111; B = 8'b10001101; // Expected: {'P': 21291}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010111; B = 8'b10001101; | Outputs: P=%b | Expected: P=%d",
                 2224,
                 
                 P
                 , 
                 
                 21291
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001101; B = 8'b11100011; // Expected: {'P': 32007}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001101; B = 8'b11100011; | Outputs: P=%b | Expected: P=%d",
                 2225,
                 
                 P
                 , 
                 
                 32007
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100100; B = 8'b00111100; // Expected: {'P': 6000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100100; B = 8'b00111100; | Outputs: P=%b | Expected: P=%d",
                 2226,
                 
                 P
                 , 
                 
                 6000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111100; B = 8'b01011101; // Expected: {'P': 11532}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111100; B = 8'b01011101; | Outputs: P=%b | Expected: P=%d",
                 2227,
                 
                 P
                 , 
                 
                 11532
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100100; B = 8'b11011001; // Expected: {'P': 35588}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100100; B = 8'b11011001; | Outputs: P=%b | Expected: P=%d",
                 2228,
                 
                 P
                 , 
                 
                 35588
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111010; B = 8'b11000110; // Expected: {'P': 36828}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111010; B = 8'b11000110; | Outputs: P=%b | Expected: P=%d",
                 2229,
                 
                 P
                 , 
                 
                 36828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100000; B = 8'b01010101; // Expected: {'P': 8160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100000; B = 8'b01010101; | Outputs: P=%b | Expected: P=%d",
                 2230,
                 
                 P
                 , 
                 
                 8160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110101; B = 8'b11111110; // Expected: {'P': 13462}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110101; B = 8'b11111110; | Outputs: P=%b | Expected: P=%d",
                 2231,
                 
                 P
                 , 
                 
                 13462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101011; B = 8'b11101011; // Expected: {'P': 10105}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101011; B = 8'b11101011; | Outputs: P=%b | Expected: P=%d",
                 2232,
                 
                 P
                 , 
                 
                 10105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110111; B = 8'b01101101; // Expected: {'P': 26923}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110111; B = 8'b01101101; | Outputs: P=%b | Expected: P=%d",
                 2233,
                 
                 P
                 , 
                 
                 26923
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100011; B = 8'b00100010; // Expected: {'P': 7718}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100011; B = 8'b00100010; | Outputs: P=%b | Expected: P=%d",
                 2234,
                 
                 P
                 , 
                 
                 7718
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101100; B = 8'b01010101; // Expected: {'P': 3740}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101100; B = 8'b01010101; | Outputs: P=%b | Expected: P=%d",
                 2235,
                 
                 P
                 , 
                 
                 3740
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001000; B = 8'b10010110; // Expected: {'P': 30000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001000; B = 8'b10010110; | Outputs: P=%b | Expected: P=%d",
                 2236,
                 
                 P
                 , 
                 
                 30000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111001; B = 8'b10000000; // Expected: {'P': 31872}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111001; B = 8'b10000000; | Outputs: P=%b | Expected: P=%d",
                 2237,
                 
                 P
                 , 
                 
                 31872
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000111; B = 8'b01011111; // Expected: {'P': 665}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000111; B = 8'b01011111; | Outputs: P=%b | Expected: P=%d",
                 2238,
                 
                 P
                 , 
                 
                 665
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110110; B = 8'b00101011; // Expected: {'P': 2322}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110110; B = 8'b00101011; | Outputs: P=%b | Expected: P=%d",
                 2239,
                 
                 P
                 , 
                 
                 2322
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110001; B = 8'b10001111; // Expected: {'P': 34463}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110001; B = 8'b10001111; | Outputs: P=%b | Expected: P=%d",
                 2240,
                 
                 P
                 , 
                 
                 34463
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100000; B = 8'b01100110; // Expected: {'P': 22848}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100000; B = 8'b01100110; | Outputs: P=%b | Expected: P=%d",
                 2241,
                 
                 P
                 , 
                 
                 22848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001111; B = 8'b10000011; // Expected: {'P': 10349}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001111; B = 8'b10000011; | Outputs: P=%b | Expected: P=%d",
                 2242,
                 
                 P
                 , 
                 
                 10349
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001111; B = 8'b00011010; // Expected: {'P': 5382}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001111; B = 8'b00011010; | Outputs: P=%b | Expected: P=%d",
                 2243,
                 
                 P
                 , 
                 
                 5382
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101101; B = 8'b10011000; // Expected: {'P': 6840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101101; B = 8'b10011000; | Outputs: P=%b | Expected: P=%d",
                 2244,
                 
                 P
                 , 
                 
                 6840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111101; B = 8'b11001010; // Expected: {'P': 25250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111101; B = 8'b11001010; | Outputs: P=%b | Expected: P=%d",
                 2245,
                 
                 P
                 , 
                 
                 25250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001001; B = 8'b11110000; // Expected: {'P': 17520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001001; B = 8'b11110000; | Outputs: P=%b | Expected: P=%d",
                 2246,
                 
                 P
                 , 
                 
                 17520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110100; B = 8'b00111000; // Expected: {'P': 10080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110100; B = 8'b00111000; | Outputs: P=%b | Expected: P=%d",
                 2247,
                 
                 P
                 , 
                 
                 10080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110111; B = 8'b00110011; // Expected: {'P': 2805}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110111; B = 8'b00110011; | Outputs: P=%b | Expected: P=%d",
                 2248,
                 
                 P
                 , 
                 
                 2805
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100111; B = 8'b10010100; // Expected: {'P': 24716}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100111; B = 8'b10010100; | Outputs: P=%b | Expected: P=%d",
                 2249,
                 
                 P
                 , 
                 
                 24716
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000010; B = 8'b01001010; // Expected: {'P': 148}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000010; B = 8'b01001010; | Outputs: P=%b | Expected: P=%d",
                 2250,
                 
                 P
                 , 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111111; B = 8'b01111010; // Expected: {'P': 7686}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111111; B = 8'b01111010; | Outputs: P=%b | Expected: P=%d",
                 2251,
                 
                 P
                 , 
                 
                 7686
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111000; B = 8'b00010000; // Expected: {'P': 2944}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111000; B = 8'b00010000; | Outputs: P=%b | Expected: P=%d",
                 2252,
                 
                 P
                 , 
                 
                 2944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001000; B = 8'b00000100; // Expected: {'P': 800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001000; B = 8'b00000100; | Outputs: P=%b | Expected: P=%d",
                 2253,
                 
                 P
                 , 
                 
                 800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001101; B = 8'b00111100; // Expected: {'P': 12300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001101; B = 8'b00111100; | Outputs: P=%b | Expected: P=%d",
                 2254,
                 
                 P
                 , 
                 
                 12300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000110; B = 8'b00111010; // Expected: {'P': 7772}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000110; B = 8'b00111010; | Outputs: P=%b | Expected: P=%d",
                 2255,
                 
                 P
                 , 
                 
                 7772
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001110; B = 8'b00011100; // Expected: {'P': 392}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001110; B = 8'b00011100; | Outputs: P=%b | Expected: P=%d",
                 2256,
                 
                 P
                 , 
                 
                 392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111010; B = 8'b10001001; // Expected: {'P': 16714}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111010; B = 8'b10001001; | Outputs: P=%b | Expected: P=%d",
                 2257,
                 
                 P
                 , 
                 
                 16714
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000101; B = 8'b11011101; // Expected: {'P': 43537}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000101; B = 8'b11011101; | Outputs: P=%b | Expected: P=%d",
                 2258,
                 
                 P
                 , 
                 
                 43537
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010000; B = 8'b01100101; // Expected: {'P': 14544}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010000; B = 8'b01100101; | Outputs: P=%b | Expected: P=%d",
                 2259,
                 
                 P
                 , 
                 
                 14544
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101111; B = 8'b10011010; // Expected: {'P': 26950}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101111; B = 8'b10011010; | Outputs: P=%b | Expected: P=%d",
                 2260,
                 
                 P
                 , 
                 
                 26950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111111; B = 8'b00000110; // Expected: {'P': 762}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111111; B = 8'b00000110; | Outputs: P=%b | Expected: P=%d",
                 2261,
                 
                 P
                 , 
                 
                 762
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111111; B = 8'b11110100; // Expected: {'P': 15372}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111111; B = 8'b11110100; | Outputs: P=%b | Expected: P=%d",
                 2262,
                 
                 P
                 , 
                 
                 15372
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001011; B = 8'b01101010; // Expected: {'P': 1166}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001011; B = 8'b01101010; | Outputs: P=%b | Expected: P=%d",
                 2263,
                 
                 P
                 , 
                 
                 1166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111100; B = 8'b00111001; // Expected: {'P': 14364}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111100; B = 8'b00111001; | Outputs: P=%b | Expected: P=%d",
                 2264,
                 
                 P
                 , 
                 
                 14364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001011; B = 8'b00001111; // Expected: {'P': 165}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001011; B = 8'b00001111; | Outputs: P=%b | Expected: P=%d",
                 2265,
                 
                 P
                 , 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001100; B = 8'b00010000; // Expected: {'P': 3264}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001100; B = 8'b00010000; | Outputs: P=%b | Expected: P=%d",
                 2266,
                 
                 P
                 , 
                 
                 3264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100001; B = 8'b11111110; // Expected: {'P': 57150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100001; B = 8'b11111110; | Outputs: P=%b | Expected: P=%d",
                 2267,
                 
                 P
                 , 
                 
                 57150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101110; B = 8'b11001110; // Expected: {'P': 22660}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101110; B = 8'b11001110; | Outputs: P=%b | Expected: P=%d",
                 2268,
                 
                 P
                 , 
                 
                 22660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100101; B = 8'b01001111; // Expected: {'P': 2923}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100101; B = 8'b01001111; | Outputs: P=%b | Expected: P=%d",
                 2269,
                 
                 P
                 , 
                 
                 2923
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110100; B = 8'b01100101; // Expected: {'P': 24644}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110100; B = 8'b01100101; | Outputs: P=%b | Expected: P=%d",
                 2270,
                 
                 P
                 , 
                 
                 24644
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110110; B = 8'b11011100; // Expected: {'P': 40040}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110110; B = 8'b11011100; | Outputs: P=%b | Expected: P=%d",
                 2271,
                 
                 P
                 , 
                 
                 40040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100000; B = 8'b11110011; // Expected: {'P': 54432}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100000; B = 8'b11110011; | Outputs: P=%b | Expected: P=%d",
                 2272,
                 
                 P
                 , 
                 
                 54432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100110; B = 8'b11011100; // Expected: {'P': 36520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100110; B = 8'b11011100; | Outputs: P=%b | Expected: P=%d",
                 2273,
                 
                 P
                 , 
                 
                 36520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001111; B = 8'b00111011; // Expected: {'P': 8437}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001111; B = 8'b00111011; | Outputs: P=%b | Expected: P=%d",
                 2274,
                 
                 P
                 , 
                 
                 8437
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001111; B = 8'b01101010; // Expected: {'P': 15158}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001111; B = 8'b01101010; | Outputs: P=%b | Expected: P=%d",
                 2275,
                 
                 P
                 , 
                 
                 15158
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010111; B = 8'b01100101; // Expected: {'P': 21715}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010111; B = 8'b01100101; | Outputs: P=%b | Expected: P=%d",
                 2276,
                 
                 P
                 , 
                 
                 21715
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010000; B = 8'b01000110; // Expected: {'P': 14560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010000; B = 8'b01000110; | Outputs: P=%b | Expected: P=%d",
                 2277,
                 
                 P
                 , 
                 
                 14560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001010; B = 8'b11111101; // Expected: {'P': 34914}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001010; B = 8'b11111101; | Outputs: P=%b | Expected: P=%d",
                 2278,
                 
                 P
                 , 
                 
                 34914
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001100; B = 8'b01011100; // Expected: {'P': 12880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001100; B = 8'b01011100; | Outputs: P=%b | Expected: P=%d",
                 2279,
                 
                 P
                 , 
                 
                 12880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111101; B = 8'b00001010; // Expected: {'P': 610}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111101; B = 8'b00001010; | Outputs: P=%b | Expected: P=%d",
                 2280,
                 
                 P
                 , 
                 
                 610
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110110; B = 8'b00010111; // Expected: {'P': 4186}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110110; B = 8'b00010111; | Outputs: P=%b | Expected: P=%d",
                 2281,
                 
                 P
                 , 
                 
                 4186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011110; B = 8'b10100100; // Expected: {'P': 15416}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011110; B = 8'b10100100; | Outputs: P=%b | Expected: P=%d",
                 2282,
                 
                 P
                 , 
                 
                 15416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000011; B = 8'b11010001; // Expected: {'P': 27379}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000011; B = 8'b11010001; | Outputs: P=%b | Expected: P=%d",
                 2283,
                 
                 P
                 , 
                 
                 27379
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100111; B = 8'b11011011; // Expected: {'P': 50589}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100111; B = 8'b11011011; | Outputs: P=%b | Expected: P=%d",
                 2284,
                 
                 P
                 , 
                 
                 50589
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101101; B = 8'b01100001; // Expected: {'P': 10573}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101101; B = 8'b01100001; | Outputs: P=%b | Expected: P=%d",
                 2285,
                 
                 P
                 , 
                 
                 10573
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011100; B = 8'b10001010; // Expected: {'P': 3864}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011100; B = 8'b10001010; | Outputs: P=%b | Expected: P=%d",
                 2286,
                 
                 P
                 , 
                 
                 3864
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100000; B = 8'b10011011; // Expected: {'P': 34720}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100000; B = 8'b10011011; | Outputs: P=%b | Expected: P=%d",
                 2287,
                 
                 P
                 , 
                 
                 34720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100110; B = 8'b00010101; // Expected: {'P': 798}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100110; B = 8'b00010101; | Outputs: P=%b | Expected: P=%d",
                 2288,
                 
                 P
                 , 
                 
                 798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111111; B = 8'b10000110; // Expected: {'P': 34170}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111111; B = 8'b10000110; | Outputs: P=%b | Expected: P=%d",
                 2289,
                 
                 P
                 , 
                 
                 34170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110111; B = 8'b00010001; // Expected: {'P': 4199}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110111; B = 8'b00010001; | Outputs: P=%b | Expected: P=%d",
                 2290,
                 
                 P
                 , 
                 
                 4199
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001001; B = 8'b00011101; // Expected: {'P': 3973}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001001; B = 8'b00011101; | Outputs: P=%b | Expected: P=%d",
                 2291,
                 
                 P
                 , 
                 
                 3973
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101110; B = 8'b11001100; // Expected: {'P': 35496}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101110; B = 8'b11001100; | Outputs: P=%b | Expected: P=%d",
                 2292,
                 
                 P
                 , 
                 
                 35496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010100; B = 8'b11001101; // Expected: {'P': 17220}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010100; B = 8'b11001101; | Outputs: P=%b | Expected: P=%d",
                 2293,
                 
                 P
                 , 
                 
                 17220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110101; B = 8'b10110010; // Expected: {'P': 9434}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110101; B = 8'b10110010; | Outputs: P=%b | Expected: P=%d",
                 2294,
                 
                 P
                 , 
                 
                 9434
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011010; B = 8'b11101010; // Expected: {'P': 51012}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011010; B = 8'b11101010; | Outputs: P=%b | Expected: P=%d",
                 2295,
                 
                 P
                 , 
                 
                 51012
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001010; B = 8'b01101001; // Expected: {'P': 1050}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001010; B = 8'b01101001; | Outputs: P=%b | Expected: P=%d",
                 2296,
                 
                 P
                 , 
                 
                 1050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001111; B = 8'b00000011; // Expected: {'P': 621}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001111; B = 8'b00000011; | Outputs: P=%b | Expected: P=%d",
                 2297,
                 
                 P
                 , 
                 
                 621
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111011; B = 8'b11110001; // Expected: {'P': 45067}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111011; B = 8'b11110001; | Outputs: P=%b | Expected: P=%d",
                 2298,
                 
                 P
                 , 
                 
                 45067
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001101; B = 8'b01000001; // Expected: {'P': 5005}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001101; B = 8'b01000001; | Outputs: P=%b | Expected: P=%d",
                 2299,
                 
                 P
                 , 
                 
                 5005
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000101; B = 8'b10011110; // Expected: {'P': 31126}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000101; B = 8'b10011110; | Outputs: P=%b | Expected: P=%d",
                 2300,
                 
                 P
                 , 
                 
                 31126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001011; B = 8'b11101011; // Expected: {'P': 2585}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001011; B = 8'b11101011; | Outputs: P=%b | Expected: P=%d",
                 2301,
                 
                 P
                 , 
                 
                 2585
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100011; B = 8'b01110001; // Expected: {'P': 25651}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100011; B = 8'b01110001; | Outputs: P=%b | Expected: P=%d",
                 2302,
                 
                 P
                 , 
                 
                 25651
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011000; B = 8'b11100011; // Expected: {'P': 34504}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011000; B = 8'b11100011; | Outputs: P=%b | Expected: P=%d",
                 2303,
                 
                 P
                 , 
                 
                 34504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000100; B = 8'b11100110; // Expected: {'P': 30360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000100; B = 8'b11100110; | Outputs: P=%b | Expected: P=%d",
                 2304,
                 
                 P
                 , 
                 
                 30360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100101; B = 8'b11001011; // Expected: {'P': 20503}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100101; B = 8'b11001011; | Outputs: P=%b | Expected: P=%d",
                 2305,
                 
                 P
                 , 
                 
                 20503
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111011; B = 8'b11011001; // Expected: {'P': 54467}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111011; B = 8'b11011001; | Outputs: P=%b | Expected: P=%d",
                 2306,
                 
                 P
                 , 
                 
                 54467
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111111; B = 8'b01000110; // Expected: {'P': 13370}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111111; B = 8'b01000110; | Outputs: P=%b | Expected: P=%d",
                 2307,
                 
                 P
                 , 
                 
                 13370
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011111; B = 8'b10001000; // Expected: {'P': 4216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011111; B = 8'b10001000; | Outputs: P=%b | Expected: P=%d",
                 2308,
                 
                 P
                 , 
                 
                 4216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111110; B = 8'b11010000; // Expected: {'P': 12896}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111110; B = 8'b11010000; | Outputs: P=%b | Expected: P=%d",
                 2309,
                 
                 P
                 , 
                 
                 12896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011010; B = 8'b01010001; // Expected: {'P': 7290}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011010; B = 8'b01010001; | Outputs: P=%b | Expected: P=%d",
                 2310,
                 
                 P
                 , 
                 
                 7290
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000000; B = 8'b10011100; // Expected: {'P': 9984}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000000; B = 8'b10011100; | Outputs: P=%b | Expected: P=%d",
                 2311,
                 
                 P
                 , 
                 
                 9984
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110000; B = 8'b11011000; // Expected: {'P': 10368}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110000; B = 8'b11011000; | Outputs: P=%b | Expected: P=%d",
                 2312,
                 
                 P
                 , 
                 
                 10368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111101; B = 8'b10010001; // Expected: {'P': 8845}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111101; B = 8'b10010001; | Outputs: P=%b | Expected: P=%d",
                 2313,
                 
                 P
                 , 
                 
                 8845
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010010; B = 8'b00100001; // Expected: {'P': 6930}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010010; B = 8'b00100001; | Outputs: P=%b | Expected: P=%d",
                 2314,
                 
                 P
                 , 
                 
                 6930
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001101; B = 8'b00000011; // Expected: {'P': 231}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001101; B = 8'b00000011; | Outputs: P=%b | Expected: P=%d",
                 2315,
                 
                 P
                 , 
                 
                 231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110011; B = 8'b10100100; // Expected: {'P': 8364}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110011; B = 8'b10100100; | Outputs: P=%b | Expected: P=%d",
                 2316,
                 
                 P
                 , 
                 
                 8364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111110; B = 8'b00100100; // Expected: {'P': 4536}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111110; B = 8'b00100100; | Outputs: P=%b | Expected: P=%d",
                 2317,
                 
                 P
                 , 
                 
                 4536
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111001; B = 8'b11110000; // Expected: {'P': 44400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111001; B = 8'b11110000; | Outputs: P=%b | Expected: P=%d",
                 2318,
                 
                 P
                 , 
                 
                 44400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011100; B = 8'b01001000; // Expected: {'P': 15840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011100; B = 8'b01001000; | Outputs: P=%b | Expected: P=%d",
                 2319,
                 
                 P
                 , 
                 
                 15840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111000; B = 8'b01000001; // Expected: {'P': 16120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111000; B = 8'b01000001; | Outputs: P=%b | Expected: P=%d",
                 2320,
                 
                 P
                 , 
                 
                 16120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100010; B = 8'b11010110; // Expected: {'P': 20972}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100010; B = 8'b11010110; | Outputs: P=%b | Expected: P=%d",
                 2321,
                 
                 P
                 , 
                 
                 20972
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101000; B = 8'b00011100; // Expected: {'P': 6496}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101000; B = 8'b00011100; | Outputs: P=%b | Expected: P=%d",
                 2322,
                 
                 P
                 , 
                 
                 6496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001100; B = 8'b11111100; // Expected: {'P': 51408}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001100; B = 8'b11111100; | Outputs: P=%b | Expected: P=%d",
                 2323,
                 
                 P
                 , 
                 
                 51408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010100; B = 8'b01011010; // Expected: {'P': 13320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010100; B = 8'b01011010; | Outputs: P=%b | Expected: P=%d",
                 2324,
                 
                 P
                 , 
                 
                 13320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010000; B = 8'b01110000; // Expected: {'P': 23296}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010000; B = 8'b01110000; | Outputs: P=%b | Expected: P=%d",
                 2325,
                 
                 P
                 , 
                 
                 23296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101010; B = 8'b11100001; // Expected: {'P': 38250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101010; B = 8'b11100001; | Outputs: P=%b | Expected: P=%d",
                 2326,
                 
                 P
                 , 
                 
                 38250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110011; B = 8'b11001110; // Expected: {'P': 23690}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110011; B = 8'b11001110; | Outputs: P=%b | Expected: P=%d",
                 2327,
                 
                 P
                 , 
                 
                 23690
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011000; B = 8'b01011010; // Expected: {'P': 13680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011000; B = 8'b01011010; | Outputs: P=%b | Expected: P=%d",
                 2328,
                 
                 P
                 , 
                 
                 13680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010001; B = 8'b10101001; // Expected: {'P': 13689}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010001; B = 8'b10101001; | Outputs: P=%b | Expected: P=%d",
                 2329,
                 
                 P
                 , 
                 
                 13689
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110111; B = 8'b10110010; // Expected: {'P': 9790}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110111; B = 8'b10110010; | Outputs: P=%b | Expected: P=%d",
                 2330,
                 
                 P
                 , 
                 
                 9790
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110110; B = 8'b00111010; // Expected: {'P': 14268}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110110; B = 8'b00111010; | Outputs: P=%b | Expected: P=%d",
                 2331,
                 
                 P
                 , 
                 
                 14268
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001101; B = 8'b10110010; // Expected: {'P': 13706}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001101; B = 8'b10110010; | Outputs: P=%b | Expected: P=%d",
                 2332,
                 
                 P
                 , 
                 
                 13706
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101110; B = 8'b00000111; // Expected: {'P': 1666}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101110; B = 8'b00000111; | Outputs: P=%b | Expected: P=%d",
                 2333,
                 
                 P
                 , 
                 
                 1666
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100000; B = 8'b00101011; // Expected: {'P': 4128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100000; B = 8'b00101011; | Outputs: P=%b | Expected: P=%d",
                 2334,
                 
                 P
                 , 
                 
                 4128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000111; B = 8'b01001100; // Expected: {'P': 15124}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000111; B = 8'b01001100; | Outputs: P=%b | Expected: P=%d",
                 2335,
                 
                 P
                 , 
                 
                 15124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000111; B = 8'b10001001; // Expected: {'P': 959}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000111; B = 8'b10001001; | Outputs: P=%b | Expected: P=%d",
                 2336,
                 
                 P
                 , 
                 
                 959
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111100; B = 8'b01000101; // Expected: {'P': 4140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111100; B = 8'b01000101; | Outputs: P=%b | Expected: P=%d",
                 2337,
                 
                 P
                 , 
                 
                 4140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111111; B = 8'b00010110; // Expected: {'P': 2794}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111111; B = 8'b00010110; | Outputs: P=%b | Expected: P=%d",
                 2338,
                 
                 P
                 , 
                 
                 2794
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111000; B = 8'b10110010; // Expected: {'P': 32752}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111000; B = 8'b10110010; | Outputs: P=%b | Expected: P=%d",
                 2339,
                 
                 P
                 , 
                 
                 32752
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101110; B = 8'b10010100; // Expected: {'P': 16280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101110; B = 8'b10010100; | Outputs: P=%b | Expected: P=%d",
                 2340,
                 
                 P
                 , 
                 
                 16280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100100; B = 8'b00011111; // Expected: {'P': 5084}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100100; B = 8'b00011111; | Outputs: P=%b | Expected: P=%d",
                 2341,
                 
                 P
                 , 
                 
                 5084
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111001; B = 8'b01101110; // Expected: {'P': 13310}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111001; B = 8'b01101110; | Outputs: P=%b | Expected: P=%d",
                 2342,
                 
                 P
                 , 
                 
                 13310
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100011; B = 8'b10111011; // Expected: {'P': 6545}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100011; B = 8'b10111011; | Outputs: P=%b | Expected: P=%d",
                 2343,
                 
                 P
                 , 
                 
                 6545
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110101; B = 8'b01100010; // Expected: {'P': 5194}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110101; B = 8'b01100010; | Outputs: P=%b | Expected: P=%d",
                 2344,
                 
                 P
                 , 
                 
                 5194
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010110; B = 8'b10111110; // Expected: {'P': 40660}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010110; B = 8'b10111110; | Outputs: P=%b | Expected: P=%d",
                 2345,
                 
                 P
                 , 
                 
                 40660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000101; B = 8'b01100010; // Expected: {'P': 19306}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000101; B = 8'b01100010; | Outputs: P=%b | Expected: P=%d",
                 2346,
                 
                 P
                 , 
                 
                 19306
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110101; B = 8'b11010001; // Expected: {'P': 24453}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110101; B = 8'b11010001; | Outputs: P=%b | Expected: P=%d",
                 2347,
                 
                 P
                 , 
                 
                 24453
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000010; B = 8'b10101001; // Expected: {'P': 21970}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000010; B = 8'b10101001; | Outputs: P=%b | Expected: P=%d",
                 2348,
                 
                 P
                 , 
                 
                 21970
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100100; B = 8'b11101010; // Expected: {'P': 8424}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100100; B = 8'b11101010; | Outputs: P=%b | Expected: P=%d",
                 2349,
                 
                 P
                 , 
                 
                 8424
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000010; B = 8'b10101000; // Expected: {'P': 336}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000010; B = 8'b10101000; | Outputs: P=%b | Expected: P=%d",
                 2350,
                 
                 P
                 , 
                 
                 336
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101100; B = 8'b01111010; // Expected: {'P': 28792}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101100; B = 8'b01111010; | Outputs: P=%b | Expected: P=%d",
                 2351,
                 
                 P
                 , 
                 
                 28792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110010; B = 8'b11100011; // Expected: {'P': 54934}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110010; B = 8'b11100011; | Outputs: P=%b | Expected: P=%d",
                 2352,
                 
                 P
                 , 
                 
                 54934
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011001; B = 8'b00000011; // Expected: {'P': 267}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011001; B = 8'b00000011; | Outputs: P=%b | Expected: P=%d",
                 2353,
                 
                 P
                 , 
                 
                 267
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110010; B = 8'b11111111; // Expected: {'P': 29070}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110010; B = 8'b11111111; | Outputs: P=%b | Expected: P=%d",
                 2354,
                 
                 P
                 , 
                 
                 29070
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100111; B = 8'b01001001; // Expected: {'P': 2847}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100111; B = 8'b01001001; | Outputs: P=%b | Expected: P=%d",
                 2355,
                 
                 P
                 , 
                 
                 2847
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101110; B = 8'b00100110; // Expected: {'P': 9044}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101110; B = 8'b00100110; | Outputs: P=%b | Expected: P=%d",
                 2356,
                 
                 P
                 , 
                 
                 9044
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000110; B = 8'b10001010; // Expected: {'P': 828}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000110; B = 8'b10001010; | Outputs: P=%b | Expected: P=%d",
                 2357,
                 
                 P
                 , 
                 
                 828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110100; B = 8'b10011101; // Expected: {'P': 18212}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110100; B = 8'b10011101; | Outputs: P=%b | Expected: P=%d",
                 2358,
                 
                 P
                 , 
                 
                 18212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011101; B = 8'b10100000; // Expected: {'P': 4640}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011101; B = 8'b10100000; | Outputs: P=%b | Expected: P=%d",
                 2359,
                 
                 P
                 , 
                 
                 4640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100100; B = 8'b11110100; // Expected: {'P': 55632}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100100; B = 8'b11110100; | Outputs: P=%b | Expected: P=%d",
                 2360,
                 
                 P
                 , 
                 
                 55632
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010100; B = 8'b01110101; // Expected: {'P': 24804}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010100; B = 8'b01110101; | Outputs: P=%b | Expected: P=%d",
                 2361,
                 
                 P
                 , 
                 
                 24804
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110111; B = 8'b11010011; // Expected: {'P': 25109}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110111; B = 8'b11010011; | Outputs: P=%b | Expected: P=%d",
                 2362,
                 
                 P
                 , 
                 
                 25109
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110101; B = 8'b11011111; // Expected: {'P': 40363}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110101; B = 8'b11011111; | Outputs: P=%b | Expected: P=%d",
                 2363,
                 
                 P
                 , 
                 
                 40363
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110010; B = 8'b00100101; // Expected: {'P': 1850}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110010; B = 8'b00100101; | Outputs: P=%b | Expected: P=%d",
                 2364,
                 
                 P
                 , 
                 
                 1850
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100011; B = 8'b00000101; // Expected: {'P': 1135}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100011; B = 8'b00000101; | Outputs: P=%b | Expected: P=%d",
                 2365,
                 
                 P
                 , 
                 
                 1135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000001; B = 8'b10011110; // Expected: {'P': 10270}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000001; B = 8'b10011110; | Outputs: P=%b | Expected: P=%d",
                 2366,
                 
                 P
                 , 
                 
                 10270
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111111; B = 8'b11011101; // Expected: {'P': 13923}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111111; B = 8'b11011101; | Outputs: P=%b | Expected: P=%d",
                 2367,
                 
                 P
                 , 
                 
                 13923
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110111; B = 8'b01000011; // Expected: {'P': 12261}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110111; B = 8'b01000011; | Outputs: P=%b | Expected: P=%d",
                 2368,
                 
                 P
                 , 
                 
                 12261
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110111; B = 8'b10010111; // Expected: {'P': 37297}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110111; B = 8'b10010111; | Outputs: P=%b | Expected: P=%d",
                 2369,
                 
                 P
                 , 
                 
                 37297
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000111; B = 8'b11001000; // Expected: {'P': 1400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000111; B = 8'b11001000; | Outputs: P=%b | Expected: P=%d",
                 2370,
                 
                 P
                 , 
                 
                 1400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100100; B = 8'b01110011; // Expected: {'P': 11500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100100; B = 8'b01110011; | Outputs: P=%b | Expected: P=%d",
                 2371,
                 
                 P
                 , 
                 
                 11500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110100; B = 8'b00111001; // Expected: {'P': 13908}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110100; B = 8'b00111001; | Outputs: P=%b | Expected: P=%d",
                 2372,
                 
                 P
                 , 
                 
                 13908
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110111; B = 8'b10001110; // Expected: {'P': 35074}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110111; B = 8'b10001110; | Outputs: P=%b | Expected: P=%d",
                 2373,
                 
                 P
                 , 
                 
                 35074
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111111; B = 8'b01001110; // Expected: {'P': 19890}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111111; B = 8'b01001110; | Outputs: P=%b | Expected: P=%d",
                 2374,
                 
                 P
                 , 
                 
                 19890
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111000; B = 8'b01010000; // Expected: {'P': 19840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111000; B = 8'b01010000; | Outputs: P=%b | Expected: P=%d",
                 2375,
                 
                 P
                 , 
                 
                 19840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011001; B = 8'b01000011; // Expected: {'P': 10251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011001; B = 8'b01000011; | Outputs: P=%b | Expected: P=%d",
                 2376,
                 
                 P
                 , 
                 
                 10251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101111; B = 8'b00001110; // Expected: {'P': 3346}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101111; B = 8'b00001110; | Outputs: P=%b | Expected: P=%d",
                 2377,
                 
                 P
                 , 
                 
                 3346
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010010; B = 8'b10010110; // Expected: {'P': 2700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010010; B = 8'b10010110; | Outputs: P=%b | Expected: P=%d",
                 2378,
                 
                 P
                 , 
                 
                 2700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010100; B = 8'b01101100; // Expected: {'P': 22896}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010100; B = 8'b01101100; | Outputs: P=%b | Expected: P=%d",
                 2379,
                 
                 P
                 , 
                 
                 22896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011111; B = 8'b11110011; // Expected: {'P': 23085}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011111; B = 8'b11110011; | Outputs: P=%b | Expected: P=%d",
                 2380,
                 
                 P
                 , 
                 
                 23085
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011100; B = 8'b10110110; // Expected: {'P': 40040}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011100; B = 8'b10110110; | Outputs: P=%b | Expected: P=%d",
                 2381,
                 
                 P
                 , 
                 
                 40040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111011; B = 8'b01011100; // Expected: {'P': 5428}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111011; B = 8'b01011100; | Outputs: P=%b | Expected: P=%d",
                 2382,
                 
                 P
                 , 
                 
                 5428
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011001; B = 8'b01001110; // Expected: {'P': 1950}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011001; B = 8'b01001110; | Outputs: P=%b | Expected: P=%d",
                 2383,
                 
                 P
                 , 
                 
                 1950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011110; B = 8'b01011101; // Expected: {'P': 2790}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011110; B = 8'b01011101; | Outputs: P=%b | Expected: P=%d",
                 2384,
                 
                 P
                 , 
                 
                 2790
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010111; B = 8'b01000111; // Expected: {'P': 10721}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010111; B = 8'b01000111; | Outputs: P=%b | Expected: P=%d",
                 2385,
                 
                 P
                 , 
                 
                 10721
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011011; B = 8'b10011111; // Expected: {'P': 4293}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011011; B = 8'b10011111; | Outputs: P=%b | Expected: P=%d",
                 2386,
                 
                 P
                 , 
                 
                 4293
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101110; B = 8'b10100001; // Expected: {'P': 38318}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101110; B = 8'b10100001; | Outputs: P=%b | Expected: P=%d",
                 2387,
                 
                 P
                 , 
                 
                 38318
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100011; B = 8'b10010000; // Expected: {'P': 32688}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100011; B = 8'b10010000; | Outputs: P=%b | Expected: P=%d",
                 2388,
                 
                 P
                 , 
                 
                 32688
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100010; B = 8'b00101000; // Expected: {'P': 1360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100010; B = 8'b00101000; | Outputs: P=%b | Expected: P=%d",
                 2389,
                 
                 P
                 , 
                 
                 1360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001111; B = 8'b00011110; // Expected: {'P': 2370}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001111; B = 8'b00011110; | Outputs: P=%b | Expected: P=%d",
                 2390,
                 
                 P
                 , 
                 
                 2370
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000001; B = 8'b01001000; // Expected: {'P': 13896}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000001; B = 8'b01001000; | Outputs: P=%b | Expected: P=%d",
                 2391,
                 
                 P
                 , 
                 
                 13896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010010; B = 8'b00001100; // Expected: {'P': 2520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010010; B = 8'b00001100; | Outputs: P=%b | Expected: P=%d",
                 2392,
                 
                 P
                 , 
                 
                 2520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111011; B = 8'b10100101; // Expected: {'P': 20295}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111011; B = 8'b10100101; | Outputs: P=%b | Expected: P=%d",
                 2393,
                 
                 P
                 , 
                 
                 20295
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111110; B = 8'b11110110; // Expected: {'P': 30996}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111110; B = 8'b11110110; | Outputs: P=%b | Expected: P=%d",
                 2394,
                 
                 P
                 , 
                 
                 30996
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101001; B = 8'b11110111; // Expected: {'P': 25935}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101001; B = 8'b11110111; | Outputs: P=%b | Expected: P=%d",
                 2395,
                 
                 P
                 , 
                 
                 25935
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110100; B = 8'b11000010; // Expected: {'P': 10088}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110100; B = 8'b11000010; | Outputs: P=%b | Expected: P=%d",
                 2396,
                 
                 P
                 , 
                 
                 10088
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110000; B = 8'b11001011; // Expected: {'P': 48720}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110000; B = 8'b11001011; | Outputs: P=%b | Expected: P=%d",
                 2397,
                 
                 P
                 , 
                 
                 48720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001000; B = 8'b10000111; // Expected: {'P': 18360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001000; B = 8'b10000111; | Outputs: P=%b | Expected: P=%d",
                 2398,
                 
                 P
                 , 
                 
                 18360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000001; B = 8'b10011000; // Expected: {'P': 152}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000001; B = 8'b10011000; | Outputs: P=%b | Expected: P=%d",
                 2399,
                 
                 P
                 , 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101000; B = 8'b11010101; // Expected: {'P': 8520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101000; B = 8'b11010101; | Outputs: P=%b | Expected: P=%d",
                 2400,
                 
                 P
                 , 
                 
                 8520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111010; B = 8'b11100110; // Expected: {'P': 57500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111010; B = 8'b11100110; | Outputs: P=%b | Expected: P=%d",
                 2401,
                 
                 P
                 , 
                 
                 57500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001001; B = 8'b00000101; // Expected: {'P': 1005}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001001; B = 8'b00000101; | Outputs: P=%b | Expected: P=%d",
                 2402,
                 
                 P
                 , 
                 
                 1005
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000011; B = 8'b10010100; // Expected: {'P': 28860}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000011; B = 8'b10010100; | Outputs: P=%b | Expected: P=%d",
                 2403,
                 
                 P
                 , 
                 
                 28860
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001111; B = 8'b10000101; // Expected: {'P': 1995}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001111; B = 8'b10000101; | Outputs: P=%b | Expected: P=%d",
                 2404,
                 
                 P
                 , 
                 
                 1995
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11001110; B = 8'b11011000; // Expected: {'P': 44496}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11001110; B = 8'b11011000; | Outputs: P=%b | Expected: P=%d",
                 2405,
                 
                 P
                 , 
                 
                 44496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001000; B = 8'b01111001; // Expected: {'P': 16456}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001000; B = 8'b01111001; | Outputs: P=%b | Expected: P=%d",
                 2406,
                 
                 P
                 , 
                 
                 16456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101000; B = 8'b01011000; // Expected: {'P': 3520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101000; B = 8'b01011000; | Outputs: P=%b | Expected: P=%d",
                 2407,
                 
                 P
                 , 
                 
                 3520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010110; B = 8'b10011100; // Expected: {'P': 3432}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010110; B = 8'b10011100; | Outputs: P=%b | Expected: P=%d",
                 2408,
                 
                 P
                 , 
                 
                 3432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010000; B = 8'b10100001; // Expected: {'P': 33488}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010000; B = 8'b10100001; | Outputs: P=%b | Expected: P=%d",
                 2409,
                 
                 P
                 , 
                 
                 33488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000001; B = 8'b10100101; // Expected: {'P': 10725}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000001; B = 8'b10100101; | Outputs: P=%b | Expected: P=%d",
                 2410,
                 
                 P
                 , 
                 
                 10725
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111010; B = 8'b00100010; // Expected: {'P': 8500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111010; B = 8'b00100010; | Outputs: P=%b | Expected: P=%d",
                 2411,
                 
                 P
                 , 
                 
                 8500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000000; B = 8'b11000110; // Expected: {'P': 38016}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000000; B = 8'b11000110; | Outputs: P=%b | Expected: P=%d",
                 2412,
                 
                 P
                 , 
                 
                 38016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011111; B = 8'b10000100; // Expected: {'P': 12540}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011111; B = 8'b10000100; | Outputs: P=%b | Expected: P=%d",
                 2413,
                 
                 P
                 , 
                 
                 12540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010001; B = 8'b01011110; // Expected: {'P': 7614}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010001; B = 8'b01011110; | Outputs: P=%b | Expected: P=%d",
                 2414,
                 
                 P
                 , 
                 
                 7614
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000011; B = 8'b11011000; // Expected: {'P': 28296}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000011; B = 8'b11011000; | Outputs: P=%b | Expected: P=%d",
                 2415,
                 
                 P
                 , 
                 
                 28296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101010; B = 8'b10011000; // Expected: {'P': 35568}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101010; B = 8'b10011000; | Outputs: P=%b | Expected: P=%d",
                 2416,
                 
                 P
                 , 
                 
                 35568
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100110; B = 8'b00101000; // Expected: {'P': 1520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100110; B = 8'b00101000; | Outputs: P=%b | Expected: P=%d",
                 2417,
                 
                 P
                 , 
                 
                 1520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111101; B = 8'b11111001; // Expected: {'P': 31125}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111101; B = 8'b11111001; | Outputs: P=%b | Expected: P=%d",
                 2418,
                 
                 P
                 , 
                 
                 31125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111111; B = 8'b01001100; // Expected: {'P': 19380}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111111; B = 8'b01001100; | Outputs: P=%b | Expected: P=%d",
                 2419,
                 
                 P
                 , 
                 
                 19380
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011100; B = 8'b00010011; // Expected: {'P': 1748}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011100; B = 8'b00010011; | Outputs: P=%b | Expected: P=%d",
                 2420,
                 
                 P
                 , 
                 
                 1748
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010110; B = 8'b10101000; // Expected: {'P': 25200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010110; B = 8'b10101000; | Outputs: P=%b | Expected: P=%d",
                 2421,
                 
                 P
                 , 
                 
                 25200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100010; B = 8'b10101110; // Expected: {'P': 17052}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100010; B = 8'b10101110; | Outputs: P=%b | Expected: P=%d",
                 2422,
                 
                 P
                 , 
                 
                 17052
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001101; B = 8'b01000001; // Expected: {'P': 9165}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001101; B = 8'b01000001; | Outputs: P=%b | Expected: P=%d",
                 2423,
                 
                 P
                 , 
                 
                 9165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100011; B = 8'b00110011; // Expected: {'P': 11577}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100011; B = 8'b00110011; | Outputs: P=%b | Expected: P=%d",
                 2424,
                 
                 P
                 , 
                 
                 11577
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110101; B = 8'b01100001; // Expected: {'P': 23765}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110101; B = 8'b01100001; | Outputs: P=%b | Expected: P=%d",
                 2425,
                 
                 P
                 , 
                 
                 23765
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100111; B = 8'b11000100; // Expected: {'P': 7644}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100111; B = 8'b11000100; | Outputs: P=%b | Expected: P=%d",
                 2426,
                 
                 P
                 , 
                 
                 7644
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011010; B = 8'b01101001; // Expected: {'P': 22890}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011010; B = 8'b01101001; | Outputs: P=%b | Expected: P=%d",
                 2427,
                 
                 P
                 , 
                 
                 22890
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000011; B = 8'b10101111; // Expected: {'P': 11725}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000011; B = 8'b10101111; | Outputs: P=%b | Expected: P=%d",
                 2428,
                 
                 P
                 , 
                 
                 11725
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001111; B = 8'b01011011; // Expected: {'P': 1365}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001111; B = 8'b01011011; | Outputs: P=%b | Expected: P=%d",
                 2429,
                 
                 P
                 , 
                 
                 1365
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000110; B = 8'b01100010; // Expected: {'P': 6860}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000110; B = 8'b01100010; | Outputs: P=%b | Expected: P=%d",
                 2430,
                 
                 P
                 , 
                 
                 6860
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100010; B = 8'b11111010; // Expected: {'P': 40500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100010; B = 8'b11111010; | Outputs: P=%b | Expected: P=%d",
                 2431,
                 
                 P
                 , 
                 
                 40500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010011; B = 8'b11111010; // Expected: {'P': 52750}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010011; B = 8'b11111010; | Outputs: P=%b | Expected: P=%d",
                 2432,
                 
                 P
                 , 
                 
                 52750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100000; B = 8'b00010011; // Expected: {'P': 4256}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100000; B = 8'b00010011; | Outputs: P=%b | Expected: P=%d",
                 2433,
                 
                 P
                 , 
                 
                 4256
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110101; B = 8'b11001000; // Expected: {'P': 23400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110101; B = 8'b11001000; | Outputs: P=%b | Expected: P=%d",
                 2434,
                 
                 P
                 , 
                 
                 23400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110011; B = 8'b10101000; // Expected: {'P': 30072}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110011; B = 8'b10101000; | Outputs: P=%b | Expected: P=%d",
                 2435,
                 
                 P
                 , 
                 
                 30072
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010110; B = 8'b00101101; // Expected: {'P': 990}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010110; B = 8'b00101101; | Outputs: P=%b | Expected: P=%d",
                 2436,
                 
                 P
                 , 
                 
                 990
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011001; B = 8'b01011001; // Expected: {'P': 19313}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011001; B = 8'b01011001; | Outputs: P=%b | Expected: P=%d",
                 2437,
                 
                 P
                 , 
                 
                 19313
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011110; B = 8'b00000110; // Expected: {'P': 180}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011110; B = 8'b00000110; | Outputs: P=%b | Expected: P=%d",
                 2438,
                 
                 P
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011100; B = 8'b10001011; // Expected: {'P': 12788}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011100; B = 8'b10001011; | Outputs: P=%b | Expected: P=%d",
                 2439,
                 
                 P
                 , 
                 
                 12788
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000001; B = 8'b11100011; // Expected: {'P': 43811}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000001; B = 8'b11100011; | Outputs: P=%b | Expected: P=%d",
                 2440,
                 
                 P
                 , 
                 
                 43811
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101100; B = 8'b11101101; // Expected: {'P': 25596}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101100; B = 8'b11101101; | Outputs: P=%b | Expected: P=%d",
                 2441,
                 
                 P
                 , 
                 
                 25596
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001011; B = 8'b11000101; // Expected: {'P': 27383}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001011; B = 8'b11000101; | Outputs: P=%b | Expected: P=%d",
                 2442,
                 
                 P
                 , 
                 
                 27383
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111010; B = 8'b11110000; // Expected: {'P': 44640}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111010; B = 8'b11110000; | Outputs: P=%b | Expected: P=%d",
                 2443,
                 
                 P
                 , 
                 
                 44640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111010; B = 8'b00000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111010; B = 8'b00000000; | Outputs: P=%b | Expected: P=%d",
                 2444,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111101; B = 8'b00111010; // Expected: {'P': 14674}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111101; B = 8'b00111010; | Outputs: P=%b | Expected: P=%d",
                 2445,
                 
                 P
                 , 
                 
                 14674
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110111; B = 8'b10111110; // Expected: {'P': 34770}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110111; B = 8'b10111110; | Outputs: P=%b | Expected: P=%d",
                 2446,
                 
                 P
                 , 
                 
                 34770
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110110; B = 8'b01100000; // Expected: {'P': 5184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110110; B = 8'b01100000; | Outputs: P=%b | Expected: P=%d",
                 2447,
                 
                 P
                 , 
                 
                 5184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001010; B = 8'b00010101; // Expected: {'P': 2898}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001010; B = 8'b00010101; | Outputs: P=%b | Expected: P=%d",
                 2448,
                 
                 P
                 , 
                 
                 2898
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100100; B = 8'b10110000; // Expected: {'P': 40128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100100; B = 8'b10110000; | Outputs: P=%b | Expected: P=%d",
                 2449,
                 
                 P
                 , 
                 
                 40128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110101; B = 8'b11000101; // Expected: {'P': 35657}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110101; B = 8'b11000101; | Outputs: P=%b | Expected: P=%d",
                 2450,
                 
                 P
                 , 
                 
                 35657
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100010; B = 8'b10011010; // Expected: {'P': 15092}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100010; B = 8'b10011010; | Outputs: P=%b | Expected: P=%d",
                 2451,
                 
                 P
                 , 
                 
                 15092
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101110; B = 8'b00000100; // Expected: {'P': 184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101110; B = 8'b00000100; | Outputs: P=%b | Expected: P=%d",
                 2452,
                 
                 P
                 , 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101000; B = 8'b11111011; // Expected: {'P': 58232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101000; B = 8'b11111011; | Outputs: P=%b | Expected: P=%d",
                 2453,
                 
                 P
                 , 
                 
                 58232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010101; B = 8'b01101101; // Expected: {'P': 9265}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010101; B = 8'b01101101; | Outputs: P=%b | Expected: P=%d",
                 2454,
                 
                 P
                 , 
                 
                 9265
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100010; B = 8'b11100111; // Expected: {'P': 22638}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100010; B = 8'b11100111; | Outputs: P=%b | Expected: P=%d",
                 2455,
                 
                 P
                 , 
                 
                 22638
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010011; B = 8'b00000001; // Expected: {'P': 83}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010011; B = 8'b00000001; | Outputs: P=%b | Expected: P=%d",
                 2456,
                 
                 P
                 , 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110100; B = 8'b01111001; // Expected: {'P': 6292}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110100; B = 8'b01111001; | Outputs: P=%b | Expected: P=%d",
                 2457,
                 
                 P
                 , 
                 
                 6292
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110001; B = 8'b00100110; // Expected: {'P': 1862}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110001; B = 8'b00100110; | Outputs: P=%b | Expected: P=%d",
                 2458,
                 
                 P
                 , 
                 
                 1862
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011010; B = 8'b11011010; // Expected: {'P': 19620}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011010; B = 8'b11011010; | Outputs: P=%b | Expected: P=%d",
                 2459,
                 
                 P
                 , 
                 
                 19620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001100; B = 8'b10011001; // Expected: {'P': 21420}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001100; B = 8'b10011001; | Outputs: P=%b | Expected: P=%d",
                 2460,
                 
                 P
                 , 
                 
                 21420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001110; B = 8'b10000110; // Expected: {'P': 10452}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001110; B = 8'b10000110; | Outputs: P=%b | Expected: P=%d",
                 2461,
                 
                 P
                 , 
                 
                 10452
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010000; B = 8'b11000101; // Expected: {'P': 15760}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010000; B = 8'b11000101; | Outputs: P=%b | Expected: P=%d",
                 2462,
                 
                 P
                 , 
                 
                 15760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101010; B = 8'b11011001; // Expected: {'P': 23002}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101010; B = 8'b11011001; | Outputs: P=%b | Expected: P=%d",
                 2463,
                 
                 P
                 , 
                 
                 23002
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100101; B = 8'b10111011; // Expected: {'P': 30855}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100101; B = 8'b10111011; | Outputs: P=%b | Expected: P=%d",
                 2464,
                 
                 P
                 , 
                 
                 30855
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011110; B = 8'b00011111; // Expected: {'P': 2914}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011110; B = 8'b00011111; | Outputs: P=%b | Expected: P=%d",
                 2465,
                 
                 P
                 , 
                 
                 2914
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011011; B = 8'b10000001; // Expected: {'P': 3483}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011011; B = 8'b10000001; | Outputs: P=%b | Expected: P=%d",
                 2466,
                 
                 P
                 , 
                 
                 3483
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001000; B = 8'b01001010; // Expected: {'P': 592}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001000; B = 8'b01001010; | Outputs: P=%b | Expected: P=%d",
                 2467,
                 
                 P
                 , 
                 
                 592
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010100; B = 8'b10010000; // Expected: {'P': 2880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010100; B = 8'b10010000; | Outputs: P=%b | Expected: P=%d",
                 2468,
                 
                 P
                 , 
                 
                 2880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000111; B = 8'b10000101; // Expected: {'P': 9443}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000111; B = 8'b10000101; | Outputs: P=%b | Expected: P=%d",
                 2469,
                 
                 P
                 , 
                 
                 9443
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001111; B = 8'b01011111; // Expected: {'P': 7505}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001111; B = 8'b01011111; | Outputs: P=%b | Expected: P=%d",
                 2470,
                 
                 P
                 , 
                 
                 7505
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100111; B = 8'b01101001; // Expected: {'P': 10815}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100111; B = 8'b01101001; | Outputs: P=%b | Expected: P=%d",
                 2471,
                 
                 P
                 , 
                 
                 10815
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111110; B = 8'b01010111; // Expected: {'P': 22098}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111110; B = 8'b01010111; | Outputs: P=%b | Expected: P=%d",
                 2472,
                 
                 P
                 , 
                 
                 22098
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100101; B = 8'b00110100; // Expected: {'P': 11908}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100101; B = 8'b00110100; | Outputs: P=%b | Expected: P=%d",
                 2473,
                 
                 P
                 , 
                 
                 11908
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101000; B = 8'b00111010; // Expected: {'P': 9744}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101000; B = 8'b00111010; | Outputs: P=%b | Expected: P=%d",
                 2474,
                 
                 P
                 , 
                 
                 9744
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111101; B = 8'b01110110; // Expected: {'P': 7198}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111101; B = 8'b01110110; | Outputs: P=%b | Expected: P=%d",
                 2475,
                 
                 P
                 , 
                 
                 7198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111011; B = 8'b11100110; // Expected: {'P': 43010}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111011; B = 8'b11100110; | Outputs: P=%b | Expected: P=%d",
                 2476,
                 
                 P
                 , 
                 
                 43010
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011111; B = 8'b10011011; // Expected: {'P': 24645}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011111; B = 8'b10011011; | Outputs: P=%b | Expected: P=%d",
                 2477,
                 
                 P
                 , 
                 
                 24645
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000011; B = 8'b11111010; // Expected: {'P': 32750}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000011; B = 8'b11111010; | Outputs: P=%b | Expected: P=%d",
                 2478,
                 
                 P
                 , 
                 
                 32750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010101; B = 8'b11110010; // Expected: {'P': 51546}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010101; B = 8'b11110010; | Outputs: P=%b | Expected: P=%d",
                 2479,
                 
                 P
                 , 
                 
                 51546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010110; B = 8'b00100010; // Expected: {'P': 7276}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010110; B = 8'b00100010; | Outputs: P=%b | Expected: P=%d",
                 2480,
                 
                 P
                 , 
                 
                 7276
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100010; B = 8'b11011010; // Expected: {'P': 21364}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100010; B = 8'b11011010; | Outputs: P=%b | Expected: P=%d",
                 2481,
                 
                 P
                 , 
                 
                 21364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001011; B = 8'b11001010; // Expected: {'P': 15150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001011; B = 8'b11001010; | Outputs: P=%b | Expected: P=%d",
                 2482,
                 
                 P
                 , 
                 
                 15150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111110; B = 8'b11111010; // Expected: {'P': 15500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111110; B = 8'b11111010; | Outputs: P=%b | Expected: P=%d",
                 2483,
                 
                 P
                 , 
                 
                 15500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001001; B = 8'b00000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001001; B = 8'b00000000; | Outputs: P=%b | Expected: P=%d",
                 2484,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100011; B = 8'b01010100; // Expected: {'P': 13692}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100011; B = 8'b01010100; | Outputs: P=%b | Expected: P=%d",
                 2485,
                 
                 P
                 , 
                 
                 13692
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000110; B = 8'b00010001; // Expected: {'P': 1190}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000110; B = 8'b00010001; | Outputs: P=%b | Expected: P=%d",
                 2486,
                 
                 P
                 , 
                 
                 1190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101001; B = 8'b00011011; // Expected: {'P': 6291}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101001; B = 8'b00011011; | Outputs: P=%b | Expected: P=%d",
                 2487,
                 
                 P
                 , 
                 
                 6291
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001111; B = 8'b10111101; // Expected: {'P': 14931}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001111; B = 8'b10111101; | Outputs: P=%b | Expected: P=%d",
                 2488,
                 
                 P
                 , 
                 
                 14931
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011111; B = 8'b00111111; // Expected: {'P': 14049}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011111; B = 8'b00111111; | Outputs: P=%b | Expected: P=%d",
                 2489,
                 
                 P
                 , 
                 
                 14049
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010100; B = 8'b00100011; // Expected: {'P': 2940}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010100; B = 8'b00100011; | Outputs: P=%b | Expected: P=%d",
                 2490,
                 
                 P
                 , 
                 
                 2940
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011110; B = 8'b10100001; // Expected: {'P': 25438}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011110; B = 8'b10100001; | Outputs: P=%b | Expected: P=%d",
                 2491,
                 
                 P
                 , 
                 
                 25438
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111011; B = 8'b11101000; // Expected: {'P': 13688}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111011; B = 8'b11101000; | Outputs: P=%b | Expected: P=%d",
                 2492,
                 
                 P
                 , 
                 
                 13688
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001011; B = 8'b01000011; // Expected: {'P': 737}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001011; B = 8'b01000011; | Outputs: P=%b | Expected: P=%d",
                 2493,
                 
                 P
                 , 
                 
                 737
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000100; B = 8'b10100001; // Expected: {'P': 21252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000100; B = 8'b10100001; | Outputs: P=%b | Expected: P=%d",
                 2494,
                 
                 P
                 , 
                 
                 21252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011110; B = 8'b00101110; // Expected: {'P': 10212}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011110; B = 8'b00101110; | Outputs: P=%b | Expected: P=%d",
                 2495,
                 
                 P
                 , 
                 
                 10212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110000; B = 8'b00001101; // Expected: {'P': 3120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110000; B = 8'b00001101; | Outputs: P=%b | Expected: P=%d",
                 2496,
                 
                 P
                 , 
                 
                 3120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011010; B = 8'b10110111; // Expected: {'P': 39894}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011010; B = 8'b10110111; | Outputs: P=%b | Expected: P=%d",
                 2497,
                 
                 P
                 , 
                 
                 39894
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001111; B = 8'b10001010; // Expected: {'P': 19734}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001111; B = 8'b10001010; | Outputs: P=%b | Expected: P=%d",
                 2498,
                 
                 P
                 , 
                 
                 19734
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000110; B = 8'b01010100; // Expected: {'P': 5880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000110; B = 8'b01010100; | Outputs: P=%b | Expected: P=%d",
                 2499,
                 
                 P
                 , 
                 
                 5880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101000; B = 8'b01000100; // Expected: {'P': 15776}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101000; B = 8'b01000100; | Outputs: P=%b | Expected: P=%d",
                 2500,
                 
                 P
                 , 
                 
                 15776
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111110; B = 8'b10100110; // Expected: {'P': 10292}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111110; B = 8'b10100110; | Outputs: P=%b | Expected: P=%d",
                 2501,
                 
                 P
                 , 
                 
                 10292
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101110; B = 8'b00101110; // Expected: {'P': 8004}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101110; B = 8'b00101110; | Outputs: P=%b | Expected: P=%d",
                 2502,
                 
                 P
                 , 
                 
                 8004
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101010; B = 8'b11000111; // Expected: {'P': 33830}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101010; B = 8'b11000111; | Outputs: P=%b | Expected: P=%d",
                 2503,
                 
                 P
                 , 
                 
                 33830
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011101; B = 8'b01100110; // Expected: {'P': 2958}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011101; B = 8'b01100110; | Outputs: P=%b | Expected: P=%d",
                 2504,
                 
                 P
                 , 
                 
                 2958
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011110; B = 8'b11111100; // Expected: {'P': 7560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011110; B = 8'b11111100; | Outputs: P=%b | Expected: P=%d",
                 2505,
                 
                 P
                 , 
                 
                 7560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010100; B = 8'b10011101; // Expected: {'P': 3140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010100; B = 8'b10011101; | Outputs: P=%b | Expected: P=%d",
                 2506,
                 
                 P
                 , 
                 
                 3140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101000; B = 8'b01100111; // Expected: {'P': 23896}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101000; B = 8'b01100111; | Outputs: P=%b | Expected: P=%d",
                 2507,
                 
                 P
                 , 
                 
                 23896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001110; B = 8'b10101010; // Expected: {'P': 13260}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001110; B = 8'b10101010; | Outputs: P=%b | Expected: P=%d",
                 2508,
                 
                 P
                 , 
                 
                 13260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101101; B = 8'b10100100; // Expected: {'P': 28372}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101101; B = 8'b10100100; | Outputs: P=%b | Expected: P=%d",
                 2509,
                 
                 P
                 , 
                 
                 28372
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011110; B = 8'b01001111; // Expected: {'P': 7426}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011110; B = 8'b01001111; | Outputs: P=%b | Expected: P=%d",
                 2510,
                 
                 P
                 , 
                 
                 7426
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011101; B = 8'b01010000; // Expected: {'P': 12560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011101; B = 8'b01010000; | Outputs: P=%b | Expected: P=%d",
                 2511,
                 
                 P
                 , 
                 
                 12560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010010; B = 8'b01100011; // Expected: {'P': 14454}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010010; B = 8'b01100011; | Outputs: P=%b | Expected: P=%d",
                 2512,
                 
                 P
                 , 
                 
                 14454
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011111; B = 8'b10000100; // Expected: {'P': 20988}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011111; B = 8'b10000100; | Outputs: P=%b | Expected: P=%d",
                 2513,
                 
                 P
                 , 
                 
                 20988
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111100; B = 8'b01110010; // Expected: {'P': 6840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111100; B = 8'b01110010; | Outputs: P=%b | Expected: P=%d",
                 2514,
                 
                 P
                 , 
                 
                 6840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111001; B = 8'b10101100; // Expected: {'P': 42828}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111001; B = 8'b10101100; | Outputs: P=%b | Expected: P=%d",
                 2515,
                 
                 P
                 , 
                 
                 42828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001100; B = 8'b01001001; // Expected: {'P': 10220}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001100; B = 8'b01001001; | Outputs: P=%b | Expected: P=%d",
                 2516,
                 
                 P
                 , 
                 
                 10220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110001; B = 8'b11001111; // Expected: {'P': 36639}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110001; B = 8'b11001111; | Outputs: P=%b | Expected: P=%d",
                 2517,
                 
                 P
                 , 
                 
                 36639
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010010; B = 8'b00001001; // Expected: {'P': 1890}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010010; B = 8'b00001001; | Outputs: P=%b | Expected: P=%d",
                 2518,
                 
                 P
                 , 
                 
                 1890
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110100; B = 8'b01110000; // Expected: {'P': 20160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110100; B = 8'b01110000; | Outputs: P=%b | Expected: P=%d",
                 2519,
                 
                 P
                 , 
                 
                 20160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101010; B = 8'b01100001; // Expected: {'P': 10282}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101010; B = 8'b01100001; | Outputs: P=%b | Expected: P=%d",
                 2520,
                 
                 P
                 , 
                 
                 10282
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011111; B = 8'b11010101; // Expected: {'P': 6603}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011111; B = 8'b11010101; | Outputs: P=%b | Expected: P=%d",
                 2521,
                 
                 P
                 , 
                 
                 6603
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010100; B = 8'b11010101; // Expected: {'P': 17892}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010100; B = 8'b11010101; | Outputs: P=%b | Expected: P=%d",
                 2522,
                 
                 P
                 , 
                 
                 17892
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110001; B = 8'b00001000; // Expected: {'P': 1416}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110001; B = 8'b00001000; | Outputs: P=%b | Expected: P=%d",
                 2523,
                 
                 P
                 , 
                 
                 1416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101100; B = 8'b11010001; // Expected: {'P': 9196}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101100; B = 8'b11010001; | Outputs: P=%b | Expected: P=%d",
                 2524,
                 
                 P
                 , 
                 
                 9196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101111; B = 8'b10110000; // Expected: {'P': 8272}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101111; B = 8'b10110000; | Outputs: P=%b | Expected: P=%d",
                 2525,
                 
                 P
                 , 
                 
                 8272
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100011; B = 8'b00000010; // Expected: {'P': 198}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100011; B = 8'b00000010; | Outputs: P=%b | Expected: P=%d",
                 2526,
                 
                 P
                 , 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001000; B = 8'b01010010; // Expected: {'P': 5904}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001000; B = 8'b01010010; | Outputs: P=%b | Expected: P=%d",
                 2527,
                 
                 P
                 , 
                 
                 5904
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010001; B = 8'b10011101; // Expected: {'P': 22765}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010001; B = 8'b10011101; | Outputs: P=%b | Expected: P=%d",
                 2528,
                 
                 P
                 , 
                 
                 22765
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011010; B = 8'b11101111; // Expected: {'P': 52102}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011010; B = 8'b11101111; | Outputs: P=%b | Expected: P=%d",
                 2529,
                 
                 P
                 , 
                 
                 52102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111100; B = 8'b10010000; // Expected: {'P': 17856}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111100; B = 8'b10010000; | Outputs: P=%b | Expected: P=%d",
                 2530,
                 
                 P
                 , 
                 
                 17856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101001; B = 8'b11110001; // Expected: {'P': 40729}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101001; B = 8'b11110001; | Outputs: P=%b | Expected: P=%d",
                 2531,
                 
                 P
                 , 
                 
                 40729
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101000; B = 8'b00001100; // Expected: {'P': 480}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101000; B = 8'b00001100; | Outputs: P=%b | Expected: P=%d",
                 2532,
                 
                 P
                 , 
                 
                 480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001000; B = 8'b11000010; // Expected: {'P': 1552}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001000; B = 8'b11000010; | Outputs: P=%b | Expected: P=%d",
                 2533,
                 
                 P
                 , 
                 
                 1552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101110; B = 8'b10111110; // Expected: {'P': 33060}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101110; B = 8'b10111110; | Outputs: P=%b | Expected: P=%d",
                 2534,
                 
                 P
                 , 
                 
                 33060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010010; B = 8'b11100100; // Expected: {'P': 47880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010010; B = 8'b11100100; | Outputs: P=%b | Expected: P=%d",
                 2535,
                 
                 P
                 , 
                 
                 47880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111111; B = 8'b01010100; // Expected: {'P': 5292}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111111; B = 8'b01010100; | Outputs: P=%b | Expected: P=%d",
                 2536,
                 
                 P
                 , 
                 
                 5292
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100110; B = 8'b00010111; // Expected: {'P': 3818}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100110; B = 8'b00010111; | Outputs: P=%b | Expected: P=%d",
                 2537,
                 
                 P
                 , 
                 
                 3818
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100011; B = 8'b01110011; // Expected: {'P': 11385}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100011; B = 8'b01110011; | Outputs: P=%b | Expected: P=%d",
                 2538,
                 
                 P
                 , 
                 
                 11385
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011110; B = 8'b11000101; // Expected: {'P': 5910}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011110; B = 8'b11000101; | Outputs: P=%b | Expected: P=%d",
                 2539,
                 
                 P
                 , 
                 
                 5910
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110101; B = 8'b01110111; // Expected: {'P': 13923}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110101; B = 8'b01110111; | Outputs: P=%b | Expected: P=%d",
                 2540,
                 
                 P
                 , 
                 
                 13923
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111100; B = 8'b00011011; // Expected: {'P': 6804}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111100; B = 8'b00011011; | Outputs: P=%b | Expected: P=%d",
                 2541,
                 
                 P
                 , 
                 
                 6804
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010110; B = 8'b11000110; // Expected: {'P': 4356}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010110; B = 8'b11000110; | Outputs: P=%b | Expected: P=%d",
                 2542,
                 
                 P
                 , 
                 
                 4356
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00000011; B = 8'b00010111; // Expected: {'P': 69}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00000011; B = 8'b00010111; | Outputs: P=%b | Expected: P=%d",
                 2543,
                 
                 P
                 , 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001111; B = 8'b00010010; // Expected: {'P': 1422}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001111; B = 8'b00010010; | Outputs: P=%b | Expected: P=%d",
                 2544,
                 
                 P
                 , 
                 
                 1422
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010110; B = 8'b00110110; // Expected: {'P': 4644}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010110; B = 8'b00110110; | Outputs: P=%b | Expected: P=%d",
                 2545,
                 
                 P
                 , 
                 
                 4644
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001101; B = 8'b01100110; // Expected: {'P': 7854}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001101; B = 8'b01100110; | Outputs: P=%b | Expected: P=%d",
                 2546,
                 
                 P
                 , 
                 
                 7854
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110111; B = 8'b00011101; // Expected: {'P': 5307}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110111; B = 8'b00011101; | Outputs: P=%b | Expected: P=%d",
                 2547,
                 
                 P
                 , 
                 
                 5307
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010011; B = 8'b11100101; // Expected: {'P': 4351}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010011; B = 8'b11100101; | Outputs: P=%b | Expected: P=%d",
                 2548,
                 
                 P
                 , 
                 
                 4351
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111111; B = 8'b00111101; // Expected: {'P': 7747}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111111; B = 8'b00111101; | Outputs: P=%b | Expected: P=%d",
                 2549,
                 
                 P
                 , 
                 
                 7747
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100010; B = 8'b00010100; // Expected: {'P': 1960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100010; B = 8'b00010100; | Outputs: P=%b | Expected: P=%d",
                 2550,
                 
                 P
                 , 
                 
                 1960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000001; B = 8'b01101000; // Expected: {'P': 20072}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000001; B = 8'b01101000; | Outputs: P=%b | Expected: P=%d",
                 2551,
                 
                 P
                 , 
                 
                 20072
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101100; B = 8'b00010101; // Expected: {'P': 3612}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101100; B = 8'b00010101; | Outputs: P=%b | Expected: P=%d",
                 2552,
                 
                 P
                 , 
                 
                 3612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110000; B = 8'b10101111; // Expected: {'P': 42000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110000; B = 8'b10101111; | Outputs: P=%b | Expected: P=%d",
                 2553,
                 
                 P
                 , 
                 
                 42000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111100; B = 8'b11010010; // Expected: {'P': 52920}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111100; B = 8'b11010010; | Outputs: P=%b | Expected: P=%d",
                 2554,
                 
                 P
                 , 
                 
                 52920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111011; B = 8'b11110100; // Expected: {'P': 30012}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111011; B = 8'b11110100; | Outputs: P=%b | Expected: P=%d",
                 2555,
                 
                 P
                 , 
                 
                 30012
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110011; B = 8'b00111100; // Expected: {'P': 14580}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110011; B = 8'b00111100; | Outputs: P=%b | Expected: P=%d",
                 2556,
                 
                 P
                 , 
                 
                 14580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110000; B = 8'b10000001; // Expected: {'P': 22704}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110000; B = 8'b10000001; | Outputs: P=%b | Expected: P=%d",
                 2557,
                 
                 P
                 , 
                 
                 22704
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000111; B = 8'b10100010; // Expected: {'P': 21870}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000111; B = 8'b10100010; | Outputs: P=%b | Expected: P=%d",
                 2558,
                 
                 P
                 , 
                 
                 21870
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111011; B = 8'b11110111; // Expected: {'P': 46189}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111011; B = 8'b11110111; | Outputs: P=%b | Expected: P=%d",
                 2559,
                 
                 P
                 , 
                 
                 46189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00111011; B = 8'b00101000; // Expected: {'P': 2360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00111011; B = 8'b00101000; | Outputs: P=%b | Expected: P=%d",
                 2560,
                 
                 P
                 , 
                 
                 2360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000101; B = 8'b11001000; // Expected: {'P': 26600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000101; B = 8'b11001000; | Outputs: P=%b | Expected: P=%d",
                 2561,
                 
                 P
                 , 
                 
                 26600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010110; B = 8'b01000101; // Expected: {'P': 5934}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010110; B = 8'b01000101; | Outputs: P=%b | Expected: P=%d",
                 2562,
                 
                 P
                 , 
                 
                 5934
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110011; B = 8'b01010010; // Expected: {'P': 19926}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110011; B = 8'b01010010; | Outputs: P=%b | Expected: P=%d",
                 2563,
                 
                 P
                 , 
                 
                 19926
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111011; B = 8'b01011001; // Expected: {'P': 10947}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111011; B = 8'b01011001; | Outputs: P=%b | Expected: P=%d",
                 2564,
                 
                 P
                 , 
                 
                 10947
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101010; B = 8'b11100111; // Expected: {'P': 24486}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101010; B = 8'b11100111; | Outputs: P=%b | Expected: P=%d",
                 2565,
                 
                 P
                 , 
                 
                 24486
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101101; B = 8'b01101110; // Expected: {'P': 26070}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101101; B = 8'b01101110; | Outputs: P=%b | Expected: P=%d",
                 2566,
                 
                 P
                 , 
                 
                 26070
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101101; B = 8'b11100010; // Expected: {'P': 53562}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101101; B = 8'b11100010; | Outputs: P=%b | Expected: P=%d",
                 2567,
                 
                 P
                 , 
                 
                 53562
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001010; B = 8'b11000111; // Expected: {'P': 1990}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001010; B = 8'b11000111; | Outputs: P=%b | Expected: P=%d",
                 2568,
                 
                 P
                 , 
                 
                 1990
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111100; B = 8'b11000101; // Expected: {'P': 49644}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111100; B = 8'b11000101; | Outputs: P=%b | Expected: P=%d",
                 2569,
                 
                 P
                 , 
                 
                 49644
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110000; B = 8'b10101110; // Expected: {'P': 19488}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110000; B = 8'b10101110; | Outputs: P=%b | Expected: P=%d",
                 2570,
                 
                 P
                 , 
                 
                 19488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100110; B = 8'b00100111; // Expected: {'P': 3978}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100110; B = 8'b00100111; | Outputs: P=%b | Expected: P=%d",
                 2571,
                 
                 P
                 , 
                 
                 3978
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101111; B = 8'b00110010; // Expected: {'P': 5550}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101111; B = 8'b00110010; | Outputs: P=%b | Expected: P=%d",
                 2572,
                 
                 P
                 , 
                 
                 5550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000011; B = 8'b11101110; // Expected: {'P': 15946}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000011; B = 8'b11101110; | Outputs: P=%b | Expected: P=%d",
                 2573,
                 
                 P
                 , 
                 
                 15946
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110111; B = 8'b10110011; // Expected: {'P': 44213}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110111; B = 8'b10110011; | Outputs: P=%b | Expected: P=%d",
                 2574,
                 
                 P
                 , 
                 
                 44213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101111; B = 8'b00000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101111; B = 8'b00000000; | Outputs: P=%b | Expected: P=%d",
                 2575,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011001; B = 8'b10110010; // Expected: {'P': 15842}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011001; B = 8'b10110010; | Outputs: P=%b | Expected: P=%d",
                 2576,
                 
                 P
                 , 
                 
                 15842
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010110; B = 8'b10011010; // Expected: {'P': 13244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010110; B = 8'b10011010; | Outputs: P=%b | Expected: P=%d",
                 2577,
                 
                 P
                 , 
                 
                 13244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110000; B = 8'b01110001; // Expected: {'P': 19888}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110000; B = 8'b01110001; | Outputs: P=%b | Expected: P=%d",
                 2578,
                 
                 P
                 , 
                 
                 19888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110101; B = 8'b10010101; // Expected: {'P': 7897}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110101; B = 8'b10010101; | Outputs: P=%b | Expected: P=%d",
                 2579,
                 
                 P
                 , 
                 
                 7897
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101111; B = 8'b11110010; // Expected: {'P': 57838}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101111; B = 8'b11110010; | Outputs: P=%b | Expected: P=%d",
                 2580,
                 
                 P
                 , 
                 
                 57838
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011100; B = 8'b10001011; // Expected: {'P': 30580}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011100; B = 8'b10001011; | Outputs: P=%b | Expected: P=%d",
                 2581,
                 
                 P
                 , 
                 
                 30580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010011; B = 8'b01011011; // Expected: {'P': 13377}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010011; B = 8'b01011011; | Outputs: P=%b | Expected: P=%d",
                 2582,
                 
                 P
                 , 
                 
                 13377
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00100011; B = 8'b11111111; // Expected: {'P': 8925}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00100011; B = 8'b11111111; | Outputs: P=%b | Expected: P=%d",
                 2583,
                 
                 P
                 , 
                 
                 8925
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100111; B = 8'b10111010; // Expected: {'P': 42966}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100111; B = 8'b10111010; | Outputs: P=%b | Expected: P=%d",
                 2584,
                 
                 P
                 , 
                 
                 42966
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111001; B = 8'b01000111; // Expected: {'P': 17679}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111001; B = 8'b01000111; | Outputs: P=%b | Expected: P=%d",
                 2585,
                 
                 P
                 , 
                 
                 17679
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000110; B = 8'b11000100; // Expected: {'P': 13720}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000110; B = 8'b11000100; | Outputs: P=%b | Expected: P=%d",
                 2586,
                 
                 P
                 , 
                 
                 13720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100000; B = 8'b01000010; // Expected: {'P': 14784}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100000; B = 8'b01000010; | Outputs: P=%b | Expected: P=%d",
                 2587,
                 
                 P
                 , 
                 
                 14784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101100; B = 8'b11111111; // Expected: {'P': 27540}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101100; B = 8'b11111111; | Outputs: P=%b | Expected: P=%d",
                 2588,
                 
                 P
                 , 
                 
                 27540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000010; B = 8'b11100001; // Expected: {'P': 29250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000010; B = 8'b11100001; | Outputs: P=%b | Expected: P=%d",
                 2589,
                 
                 P
                 , 
                 
                 29250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011110; B = 8'b10111001; // Expected: {'P': 17390}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011110; B = 8'b10111001; | Outputs: P=%b | Expected: P=%d",
                 2590,
                 
                 P
                 , 
                 
                 17390
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111000; B = 8'b01001011; // Expected: {'P': 9000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111000; B = 8'b01001011; | Outputs: P=%b | Expected: P=%d",
                 2591,
                 
                 P
                 , 
                 
                 9000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01010110; B = 8'b10000100; // Expected: {'P': 11352}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01010110; B = 8'b10000100; | Outputs: P=%b | Expected: P=%d",
                 2592,
                 
                 P
                 , 
                 
                 11352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101010; B = 8'b01011101; // Expected: {'P': 9858}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101010; B = 8'b01011101; | Outputs: P=%b | Expected: P=%d",
                 2593,
                 
                 P
                 , 
                 
                 9858
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001001; B = 8'b10100011; // Expected: {'P': 1467}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001001; B = 8'b10100011; | Outputs: P=%b | Expected: P=%d",
                 2594,
                 
                 P
                 , 
                 
                 1467
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111101; B = 8'b01111111; // Expected: {'P': 24003}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111101; B = 8'b01111111; | Outputs: P=%b | Expected: P=%d",
                 2595,
                 
                 P
                 , 
                 
                 24003
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101100; B = 8'b00111010; // Expected: {'P': 2552}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101100; B = 8'b00111010; | Outputs: P=%b | Expected: P=%d",
                 2596,
                 
                 P
                 , 
                 
                 2552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000110; B = 8'b01110101; // Expected: {'P': 23166}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000110; B = 8'b01110101; | Outputs: P=%b | Expected: P=%d",
                 2597,
                 
                 P
                 , 
                 
                 23166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010110; B = 8'b11100101; // Expected: {'P': 49006}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010110; B = 8'b11100101; | Outputs: P=%b | Expected: P=%d",
                 2598,
                 
                 P
                 , 
                 
                 49006
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110110; B = 8'b10001111; // Expected: {'P': 7722}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110110; B = 8'b10001111; | Outputs: P=%b | Expected: P=%d",
                 2599,
                 
                 P
                 , 
                 
                 7722
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100001; B = 8'b10001101; // Expected: {'P': 13677}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100001; B = 8'b10001101; | Outputs: P=%b | Expected: P=%d",
                 2600,
                 
                 P
                 , 
                 
                 13677
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110110; B = 8'b01110111; // Expected: {'P': 6426}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110110; B = 8'b01110111; | Outputs: P=%b | Expected: P=%d",
                 2601,
                 
                 P
                 , 
                 
                 6426
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00101010; B = 8'b01111011; // Expected: {'P': 5166}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00101010; B = 8'b01111011; | Outputs: P=%b | Expected: P=%d",
                 2602,
                 
                 P
                 , 
                 
                 5166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011011; B = 8'b11111011; // Expected: {'P': 38905}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011011; B = 8'b11111011; | Outputs: P=%b | Expected: P=%d",
                 2603,
                 
                 P
                 , 
                 
                 38905
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000010; B = 8'b00110001; // Expected: {'P': 6370}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000010; B = 8'b00110001; | Outputs: P=%b | Expected: P=%d",
                 2604,
                 
                 P
                 , 
                 
                 6370
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111011; B = 8'b01101100; // Expected: {'P': 27108}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111011; B = 8'b01101100; | Outputs: P=%b | Expected: P=%d",
                 2605,
                 
                 P
                 , 
                 
                 27108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011011; B = 8'b01110010; // Expected: {'P': 10374}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011011; B = 8'b01110010; | Outputs: P=%b | Expected: P=%d",
                 2606,
                 
                 P
                 , 
                 
                 10374
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101010; B = 8'b00101010; // Expected: {'P': 9828}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101010; B = 8'b00101010; | Outputs: P=%b | Expected: P=%d",
                 2607,
                 
                 P
                 , 
                 
                 9828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011000; B = 8'b01100111; // Expected: {'P': 2472}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011000; B = 8'b01100111; | Outputs: P=%b | Expected: P=%d",
                 2608,
                 
                 P
                 , 
                 
                 2472
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011100; B = 8'b11001100; // Expected: {'P': 31824}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011100; B = 8'b11001100; | Outputs: P=%b | Expected: P=%d",
                 2609,
                 
                 P
                 , 
                 
                 31824
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111000; B = 8'b00101001; // Expected: {'P': 7544}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111000; B = 8'b00101001; | Outputs: P=%b | Expected: P=%d",
                 2610,
                 
                 P
                 , 
                 
                 7544
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000000; B = 8'b10111100; // Expected: {'P': 12032}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000000; B = 8'b10111100; | Outputs: P=%b | Expected: P=%d",
                 2611,
                 
                 P
                 , 
                 
                 12032
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011010; B = 8'b10000100; // Expected: {'P': 11880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011010; B = 8'b10000100; | Outputs: P=%b | Expected: P=%d",
                 2612,
                 
                 P
                 , 
                 
                 11880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001101; B = 8'b11100110; // Expected: {'P': 32430}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001101; B = 8'b11100110; | Outputs: P=%b | Expected: P=%d",
                 2613,
                 
                 P
                 , 
                 
                 32430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101000; B = 8'b00000110; // Expected: {'P': 1008}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101000; B = 8'b00000110; | Outputs: P=%b | Expected: P=%d",
                 2614,
                 
                 P
                 , 
                 
                 1008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10110011; B = 8'b01011010; // Expected: {'P': 16110}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10110011; B = 8'b01011010; | Outputs: P=%b | Expected: P=%d",
                 2615,
                 
                 P
                 , 
                 
                 16110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100111; B = 8'b10011010; // Expected: {'P': 35574}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100111; B = 8'b10011010; | Outputs: P=%b | Expected: P=%d",
                 2616,
                 
                 P
                 , 
                 
                 35574
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11000001; B = 8'b11010100; // Expected: {'P': 40916}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11000001; B = 8'b11010100; | Outputs: P=%b | Expected: P=%d",
                 2617,
                 
                 P
                 , 
                 
                 40916
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10011111; B = 8'b11000110; // Expected: {'P': 31482}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10011111; B = 8'b11000110; | Outputs: P=%b | Expected: P=%d",
                 2618,
                 
                 P
                 , 
                 
                 31482
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111010; B = 8'b00001001; // Expected: {'P': 2250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111010; B = 8'b00001001; | Outputs: P=%b | Expected: P=%d",
                 2619,
                 
                 P
                 , 
                 
                 2250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01100011; B = 8'b00101100; // Expected: {'P': 4356}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01100011; B = 8'b00101100; | Outputs: P=%b | Expected: P=%d",
                 2620,
                 
                 P
                 , 
                 
                 4356
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00011101; B = 8'b10101010; // Expected: {'P': 4930}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00011101; B = 8'b10101010; | Outputs: P=%b | Expected: P=%d",
                 2621,
                 
                 P
                 , 
                 
                 4930
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100110; B = 8'b00101000; // Expected: {'P': 6640}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100110; B = 8'b00101000; | Outputs: P=%b | Expected: P=%d",
                 2622,
                 
                 P
                 , 
                 
                 6640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001000; B = 8'b11100110; // Expected: {'P': 31280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001000; B = 8'b11100110; | Outputs: P=%b | Expected: P=%d",
                 2623,
                 
                 P
                 , 
                 
                 31280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10100101; B = 8'b00100000; // Expected: {'P': 5280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10100101; B = 8'b00100000; | Outputs: P=%b | Expected: P=%d",
                 2624,
                 
                 P
                 , 
                 
                 5280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110001; B = 8'b01111110; // Expected: {'P': 14238}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110001; B = 8'b01111110; | Outputs: P=%b | Expected: P=%d",
                 2625,
                 
                 P
                 , 
                 
                 14238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001100; B = 8'b10011000; // Expected: {'P': 1824}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001100; B = 8'b10011000; | Outputs: P=%b | Expected: P=%d",
                 2626,
                 
                 P
                 , 
                 
                 1824
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010010; B = 8'b01011100; // Expected: {'P': 13432}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010010; B = 8'b01011100; | Outputs: P=%b | Expected: P=%d",
                 2627,
                 
                 P
                 , 
                 
                 13432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011010; B = 8'b00100011; // Expected: {'P': 7630}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011010; B = 8'b00100011; | Outputs: P=%b | Expected: P=%d",
                 2628,
                 
                 P
                 , 
                 
                 7630
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100011; B = 8'b10001010; // Expected: {'P': 31326}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100011; B = 8'b10001010; | Outputs: P=%b | Expected: P=%d",
                 2629,
                 
                 P
                 , 
                 
                 31326
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011010; B = 8'b01111111; // Expected: {'P': 27686}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011010; B = 8'b01111111; | Outputs: P=%b | Expected: P=%d",
                 2630,
                 
                 P
                 , 
                 
                 27686
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10010010; B = 8'b01111111; // Expected: {'P': 18542}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10010010; B = 8'b01111111; | Outputs: P=%b | Expected: P=%d",
                 2631,
                 
                 P
                 , 
                 
                 18542
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11101111; B = 8'b10110110; // Expected: {'P': 43498}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11101111; B = 8'b10110110; | Outputs: P=%b | Expected: P=%d",
                 2632,
                 
                 P
                 , 
                 
                 43498
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101000; B = 8'b01100011; // Expected: {'P': 16632}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101000; B = 8'b01100011; | Outputs: P=%b | Expected: P=%d",
                 2633,
                 
                 P
                 , 
                 
                 16632
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00010100; B = 8'b00011001; // Expected: {'P': 500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00010100; B = 8'b00011001; | Outputs: P=%b | Expected: P=%d",
                 2634,
                 
                 P
                 , 
                 
                 500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00110001; B = 8'b01001001; // Expected: {'P': 3577}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00110001; B = 8'b01001001; | Outputs: P=%b | Expected: P=%d",
                 2635,
                 
                 P
                 , 
                 
                 3577
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010100; B = 8'b10100110; // Expected: {'P': 35192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010100; B = 8'b10100110; | Outputs: P=%b | Expected: P=%d",
                 2636,
                 
                 P
                 , 
                 
                 35192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111011; B = 8'b10111111; // Expected: {'P': 23493}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111011; B = 8'b10111111; | Outputs: P=%b | Expected: P=%d",
                 2637,
                 
                 P
                 , 
                 
                 23493
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01111110; B = 8'b01001010; // Expected: {'P': 9324}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01111110; B = 8'b01001010; | Outputs: P=%b | Expected: P=%d",
                 2638,
                 
                 P
                 , 
                 
                 9324
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01011010; B = 8'b11010011; // Expected: {'P': 18990}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01011010; B = 8'b11010011; | Outputs: P=%b | Expected: P=%d",
                 2639,
                 
                 P
                 , 
                 
                 18990
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100100; B = 8'b00010111; // Expected: {'P': 5244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100100; B = 8'b00010111; | Outputs: P=%b | Expected: P=%d",
                 2640,
                 
                 P
                 , 
                 
                 5244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001111; B = 8'b00001000; // Expected: {'P': 120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001111; B = 8'b00001000; | Outputs: P=%b | Expected: P=%d",
                 2641,
                 
                 P
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11100110; B = 8'b11000011; // Expected: {'P': 44850}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11100110; B = 8'b11000011; | Outputs: P=%b | Expected: P=%d",
                 2642,
                 
                 P
                 , 
                 
                 44850
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000000; B = 8'b01101101; // Expected: {'P': 13952}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000000; B = 8'b01101101; | Outputs: P=%b | Expected: P=%d",
                 2643,
                 
                 P
                 , 
                 
                 13952
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01110101; B = 8'b00111100; // Expected: {'P': 7020}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01110101; B = 8'b00111100; | Outputs: P=%b | Expected: P=%d",
                 2644,
                 
                 P
                 , 
                 
                 7020
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111010; B = 8'b10010111; // Expected: {'P': 37750}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111010; B = 8'b10010111; | Outputs: P=%b | Expected: P=%d",
                 2645,
                 
                 P
                 , 
                 
                 37750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10000110; B = 8'b10000001; // Expected: {'P': 17286}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10000110; B = 8'b10000001; | Outputs: P=%b | Expected: P=%d",
                 2646,
                 
                 P
                 , 
                 
                 17286
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101111; B = 8'b00111100; // Expected: {'P': 6660}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101111; B = 8'b00111100; | Outputs: P=%b | Expected: P=%d",
                 2647,
                 
                 P
                 , 
                 
                 6660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10111011; B = 8'b11000010; // Expected: {'P': 36278}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10111011; B = 8'b11000010; | Outputs: P=%b | Expected: P=%d",
                 2648,
                 
                 P
                 , 
                 
                 36278
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11011111; B = 8'b11111001; // Expected: {'P': 55527}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11011111; B = 8'b11111001; | Outputs: P=%b | Expected: P=%d",
                 2649,
                 
                 P
                 , 
                 
                 55527
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110010; B = 8'b11001100; // Expected: {'P': 49368}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110010; B = 8'b11001100; | Outputs: P=%b | Expected: P=%d",
                 2650,
                 
                 P
                 , 
                 
                 49368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10001011; B = 8'b01101010; // Expected: {'P': 14734}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10001011; B = 8'b01101010; | Outputs: P=%b | Expected: P=%d",
                 2651,
                 
                 P
                 , 
                 
                 14734
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11010011; B = 8'b11010101; // Expected: {'P': 44943}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11010011; B = 8'b11010101; | Outputs: P=%b | Expected: P=%d",
                 2652,
                 
                 P
                 , 
                 
                 44943
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11111100; B = 8'b11000010; // Expected: {'P': 48888}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11111100; B = 8'b11000010; | Outputs: P=%b | Expected: P=%d",
                 2653,
                 
                 P
                 , 
                 
                 48888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b11110101; B = 8'b11010111; // Expected: {'P': 52675}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b11110101; B = 8'b11010111; | Outputs: P=%b | Expected: P=%d",
                 2654,
                 
                 P
                 , 
                 
                 52675
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01001111; B = 8'b01111010; // Expected: {'P': 9638}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01001111; B = 8'b01111010; | Outputs: P=%b | Expected: P=%d",
                 2655,
                 
                 P
                 , 
                 
                 9638
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b00001101; B = 8'b01001000; // Expected: {'P': 936}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b00001101; B = 8'b01001000; | Outputs: P=%b | Expected: P=%d",
                 2656,
                 
                 P
                 , 
                 
                 936
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01000011; B = 8'b10100101; // Expected: {'P': 11055}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01000011; B = 8'b10100101; | Outputs: P=%b | Expected: P=%d",
                 2657,
                 
                 P
                 , 
                 
                 11055
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b01101000; B = 8'b11101001; // Expected: {'P': 24232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b01101000; B = 8'b11101001; | Outputs: P=%b | Expected: P=%d",
                 2658,
                 
                 P
                 , 
                 
                 24232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 8'b10101001; B = 8'b10101101; // Expected: {'P': 29237}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 8'b10101001; B = 8'b10101101; | Outputs: P=%b | Expected: P=%d",
                 2659,
                 
                 P
                 , 
                 
                 29237
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        $finish;
    end
  
endmodule